//  A testbench for alu_RESULT_tb
`timescale 1us/1ns

module alu_RESULT_tb;
    reg [15:0] A;
    reg [15:0] B;
    reg [1:0] ALUOP;
    wire [15:0] RESULT;
    wire [3:0] FLAG;

  alu alu0 (
    .A(A),
    .B(B),
    .ALUOP(ALUOP),
    .RESULT(RESULT),
    .FLAG(FLAG)
  );

    reg [49:0] patterns[0:5023];
    integer i;

    initial begin
      patterns[0] = 50'b00_0000000000000000_0000000000000000_0000000000000000;
      patterns[1] = 50'b01_0000000000000000_0000000000000000_0000000000000000;
      patterns[2] = 50'b10_0000000000000000_0000000000000000_0000000000000000;
      patterns[3] = 50'b11_0000000000000000_0000000000000000_0000000000000000;
      patterns[4] = 50'b00_0000000000000000_0000000000000001_0000000000000001;
      patterns[5] = 50'b01_0000000000000000_0000000000000001_1111111111111111;
      patterns[6] = 50'b10_0000000000000000_0000000000000001_0000000000000000;
      patterns[7] = 50'b11_0000000000000000_0000000000000001_0000000000000001;
      patterns[8] = 50'b00_0000000000000000_0000000000000010_0000000000000010;
      patterns[9] = 50'b01_0000000000000000_0000000000000010_1111111111111110;
      patterns[10] = 50'b10_0000000000000000_0000000000000010_0000000000000000;
      patterns[11] = 50'b11_0000000000000000_0000000000000010_0000000000000010;
      patterns[12] = 50'b00_0000000000000000_0000000000000011_0000000000000011;
      patterns[13] = 50'b01_0000000000000000_0000000000000011_1111111111111101;
      patterns[14] = 50'b10_0000000000000000_0000000000000011_0000000000000000;
      patterns[15] = 50'b11_0000000000000000_0000000000000011_0000000000000011;
      patterns[16] = 50'b00_0000000000000000_0000000000000100_0000000000000100;
      patterns[17] = 50'b01_0000000000000000_0000000000000100_1111111111111100;
      patterns[18] = 50'b10_0000000000000000_0000000000000100_0000000000000000;
      patterns[19] = 50'b11_0000000000000000_0000000000000100_0000000000000100;
      patterns[20] = 50'b00_0000000000000000_0000000000000101_0000000000000101;
      patterns[21] = 50'b01_0000000000000000_0000000000000101_1111111111111011;
      patterns[22] = 50'b10_0000000000000000_0000000000000101_0000000000000000;
      patterns[23] = 50'b11_0000000000000000_0000000000000101_0000000000000101;
      patterns[24] = 50'b00_0000000000000000_0000000000000110_0000000000000110;
      patterns[25] = 50'b01_0000000000000000_0000000000000110_1111111111111010;
      patterns[26] = 50'b10_0000000000000000_0000000000000110_0000000000000000;
      patterns[27] = 50'b11_0000000000000000_0000000000000110_0000000000000110;
      patterns[28] = 50'b00_0000000000000000_0000000000000111_0000000000000111;
      patterns[29] = 50'b01_0000000000000000_0000000000000111_1111111111111001;
      patterns[30] = 50'b10_0000000000000000_0000000000000111_0000000000000000;
      patterns[31] = 50'b11_0000000000000000_0000000000000111_0000000000000111;
      patterns[32] = 50'b00_0000000000000000_0000000000001000_0000000000001000;
      patterns[33] = 50'b01_0000000000000000_0000000000001000_1111111111111000;
      patterns[34] = 50'b10_0000000000000000_0000000000001000_0000000000000000;
      patterns[35] = 50'b11_0000000000000000_0000000000001000_0000000000001000;
      patterns[36] = 50'b00_0000000000000000_0000000000001001_0000000000001001;
      patterns[37] = 50'b01_0000000000000000_0000000000001001_1111111111110111;
      patterns[38] = 50'b10_0000000000000000_0000000000001001_0000000000000000;
      patterns[39] = 50'b11_0000000000000000_0000000000001001_0000000000001001;
      patterns[40] = 50'b00_0000000000000000_0000000000001010_0000000000001010;
      patterns[41] = 50'b01_0000000000000000_0000000000001010_1111111111110110;
      patterns[42] = 50'b10_0000000000000000_0000000000001010_0000000000000000;
      patterns[43] = 50'b11_0000000000000000_0000000000001010_0000000000001010;
      patterns[44] = 50'b00_0000000000000000_0000000000001011_0000000000001011;
      patterns[45] = 50'b01_0000000000000000_0000000000001011_1111111111110101;
      patterns[46] = 50'b10_0000000000000000_0000000000001011_0000000000000000;
      patterns[47] = 50'b11_0000000000000000_0000000000001011_0000000000001011;
      patterns[48] = 50'b00_0000000000000000_0000000000001100_0000000000001100;
      patterns[49] = 50'b01_0000000000000000_0000000000001100_1111111111110100;
      patterns[50] = 50'b10_0000000000000000_0000000000001100_0000000000000000;
      patterns[51] = 50'b11_0000000000000000_0000000000001100_0000000000001100;
      patterns[52] = 50'b00_0000000000000000_0000000000001101_0000000000001101;
      patterns[53] = 50'b01_0000000000000000_0000000000001101_1111111111110011;
      patterns[54] = 50'b10_0000000000000000_0000000000001101_0000000000000000;
      patterns[55] = 50'b11_0000000000000000_0000000000001101_0000000000001101;
      patterns[56] = 50'b00_0000000000000000_0000000000001110_0000000000001110;
      patterns[57] = 50'b01_0000000000000000_0000000000001110_1111111111110010;
      patterns[58] = 50'b10_0000000000000000_0000000000001110_0000000000000000;
      patterns[59] = 50'b11_0000000000000000_0000000000001110_0000000000001110;
      patterns[60] = 50'b00_0000000000000000_0000000000001111_0000000000001111;
      patterns[61] = 50'b01_0000000000000000_0000000000001111_1111111111110001;
      patterns[62] = 50'b10_0000000000000000_0000000000001111_0000000000000000;
      patterns[63] = 50'b11_0000000000000000_0000000000001111_0000000000001111;
      patterns[64] = 50'b00_0000000000000001_0000000000000000_0000000000000001;
      patterns[65] = 50'b01_0000000000000001_0000000000000000_0000000000000001;
      patterns[66] = 50'b10_0000000000000001_0000000000000000_0000000000000000;
      patterns[67] = 50'b11_0000000000000001_0000000000000000_0000000000000001;
      patterns[68] = 50'b00_0000000000000001_0000000000000001_0000000000000010;
      patterns[69] = 50'b01_0000000000000001_0000000000000001_0000000000000000;
      patterns[70] = 50'b10_0000000000000001_0000000000000001_0000000000000001;
      patterns[71] = 50'b11_0000000000000001_0000000000000001_0000000000000001;
      patterns[72] = 50'b00_0000000000000001_0000000000000010_0000000000000011;
      patterns[73] = 50'b01_0000000000000001_0000000000000010_1111111111111111;
      patterns[74] = 50'b10_0000000000000001_0000000000000010_0000000000000000;
      patterns[75] = 50'b11_0000000000000001_0000000000000010_0000000000000011;
      patterns[76] = 50'b00_0000000000000001_0000000000000011_0000000000000100;
      patterns[77] = 50'b01_0000000000000001_0000000000000011_1111111111111110;
      patterns[78] = 50'b10_0000000000000001_0000000000000011_0000000000000001;
      patterns[79] = 50'b11_0000000000000001_0000000000000011_0000000000000011;
      patterns[80] = 50'b00_0000000000000001_0000000000000100_0000000000000101;
      patterns[81] = 50'b01_0000000000000001_0000000000000100_1111111111111101;
      patterns[82] = 50'b10_0000000000000001_0000000000000100_0000000000000000;
      patterns[83] = 50'b11_0000000000000001_0000000000000100_0000000000000101;
      patterns[84] = 50'b00_0000000000000001_0000000000000101_0000000000000110;
      patterns[85] = 50'b01_0000000000000001_0000000000000101_1111111111111100;
      patterns[86] = 50'b10_0000000000000001_0000000000000101_0000000000000001;
      patterns[87] = 50'b11_0000000000000001_0000000000000101_0000000000000101;
      patterns[88] = 50'b00_0000000000000001_0000000000000110_0000000000000111;
      patterns[89] = 50'b01_0000000000000001_0000000000000110_1111111111111011;
      patterns[90] = 50'b10_0000000000000001_0000000000000110_0000000000000000;
      patterns[91] = 50'b11_0000000000000001_0000000000000110_0000000000000111;
      patterns[92] = 50'b00_0000000000000001_0000000000000111_0000000000001000;
      patterns[93] = 50'b01_0000000000000001_0000000000000111_1111111111111010;
      patterns[94] = 50'b10_0000000000000001_0000000000000111_0000000000000001;
      patterns[95] = 50'b11_0000000000000001_0000000000000111_0000000000000111;
      patterns[96] = 50'b00_0000000000000001_0000000000001000_0000000000001001;
      patterns[97] = 50'b01_0000000000000001_0000000000001000_1111111111111001;
      patterns[98] = 50'b10_0000000000000001_0000000000001000_0000000000000000;
      patterns[99] = 50'b11_0000000000000001_0000000000001000_0000000000001001;
      patterns[100] = 50'b00_0000000000000001_0000000000001001_0000000000001010;
      patterns[101] = 50'b01_0000000000000001_0000000000001001_1111111111111000;
      patterns[102] = 50'b10_0000000000000001_0000000000001001_0000000000000001;
      patterns[103] = 50'b11_0000000000000001_0000000000001001_0000000000001001;
      patterns[104] = 50'b00_0000000000000001_0000000000001010_0000000000001011;
      patterns[105] = 50'b01_0000000000000001_0000000000001010_1111111111110111;
      patterns[106] = 50'b10_0000000000000001_0000000000001010_0000000000000000;
      patterns[107] = 50'b11_0000000000000001_0000000000001010_0000000000001011;
      patterns[108] = 50'b00_0000000000000001_0000000000001011_0000000000001100;
      patterns[109] = 50'b01_0000000000000001_0000000000001011_1111111111110110;
      patterns[110] = 50'b10_0000000000000001_0000000000001011_0000000000000001;
      patterns[111] = 50'b11_0000000000000001_0000000000001011_0000000000001011;
      patterns[112] = 50'b00_0000000000000001_0000000000001100_0000000000001101;
      patterns[113] = 50'b01_0000000000000001_0000000000001100_1111111111110101;
      patterns[114] = 50'b10_0000000000000001_0000000000001100_0000000000000000;
      patterns[115] = 50'b11_0000000000000001_0000000000001100_0000000000001101;
      patterns[116] = 50'b00_0000000000000001_0000000000001101_0000000000001110;
      patterns[117] = 50'b01_0000000000000001_0000000000001101_1111111111110100;
      patterns[118] = 50'b10_0000000000000001_0000000000001101_0000000000000001;
      patterns[119] = 50'b11_0000000000000001_0000000000001101_0000000000001101;
      patterns[120] = 50'b00_0000000000000001_0000000000001110_0000000000001111;
      patterns[121] = 50'b01_0000000000000001_0000000000001110_1111111111110011;
      patterns[122] = 50'b10_0000000000000001_0000000000001110_0000000000000000;
      patterns[123] = 50'b11_0000000000000001_0000000000001110_0000000000001111;
      patterns[124] = 50'b00_0000000000000001_0000000000001111_0000000000010000;
      patterns[125] = 50'b01_0000000000000001_0000000000001111_1111111111110010;
      patterns[126] = 50'b10_0000000000000001_0000000000001111_0000000000000001;
      patterns[127] = 50'b11_0000000000000001_0000000000001111_0000000000001111;
      patterns[128] = 50'b00_0000000000000010_0000000000000000_0000000000000010;
      patterns[129] = 50'b01_0000000000000010_0000000000000000_0000000000000010;
      patterns[130] = 50'b10_0000000000000010_0000000000000000_0000000000000000;
      patterns[131] = 50'b11_0000000000000010_0000000000000000_0000000000000010;
      patterns[132] = 50'b00_0000000000000010_0000000000000001_0000000000000011;
      patterns[133] = 50'b01_0000000000000010_0000000000000001_0000000000000001;
      patterns[134] = 50'b10_0000000000000010_0000000000000001_0000000000000000;
      patterns[135] = 50'b11_0000000000000010_0000000000000001_0000000000000011;
      patterns[136] = 50'b00_0000000000000010_0000000000000010_0000000000000100;
      patterns[137] = 50'b01_0000000000000010_0000000000000010_0000000000000000;
      patterns[138] = 50'b10_0000000000000010_0000000000000010_0000000000000010;
      patterns[139] = 50'b11_0000000000000010_0000000000000010_0000000000000010;
      patterns[140] = 50'b00_0000000000000010_0000000000000011_0000000000000101;
      patterns[141] = 50'b01_0000000000000010_0000000000000011_1111111111111111;
      patterns[142] = 50'b10_0000000000000010_0000000000000011_0000000000000010;
      patterns[143] = 50'b11_0000000000000010_0000000000000011_0000000000000011;
      patterns[144] = 50'b00_0000000000000010_0000000000000100_0000000000000110;
      patterns[145] = 50'b01_0000000000000010_0000000000000100_1111111111111110;
      patterns[146] = 50'b10_0000000000000010_0000000000000100_0000000000000000;
      patterns[147] = 50'b11_0000000000000010_0000000000000100_0000000000000110;
      patterns[148] = 50'b00_0000000000000010_0000000000000101_0000000000000111;
      patterns[149] = 50'b01_0000000000000010_0000000000000101_1111111111111101;
      patterns[150] = 50'b10_0000000000000010_0000000000000101_0000000000000000;
      patterns[151] = 50'b11_0000000000000010_0000000000000101_0000000000000111;
      patterns[152] = 50'b00_0000000000000010_0000000000000110_0000000000001000;
      patterns[153] = 50'b01_0000000000000010_0000000000000110_1111111111111100;
      patterns[154] = 50'b10_0000000000000010_0000000000000110_0000000000000010;
      patterns[155] = 50'b11_0000000000000010_0000000000000110_0000000000000110;
      patterns[156] = 50'b00_0000000000000010_0000000000000111_0000000000001001;
      patterns[157] = 50'b01_0000000000000010_0000000000000111_1111111111111011;
      patterns[158] = 50'b10_0000000000000010_0000000000000111_0000000000000010;
      patterns[159] = 50'b11_0000000000000010_0000000000000111_0000000000000111;
      patterns[160] = 50'b00_0000000000000010_0000000000001000_0000000000001010;
      patterns[161] = 50'b01_0000000000000010_0000000000001000_1111111111111010;
      patterns[162] = 50'b10_0000000000000010_0000000000001000_0000000000000000;
      patterns[163] = 50'b11_0000000000000010_0000000000001000_0000000000001010;
      patterns[164] = 50'b00_0000000000000010_0000000000001001_0000000000001011;
      patterns[165] = 50'b01_0000000000000010_0000000000001001_1111111111111001;
      patterns[166] = 50'b10_0000000000000010_0000000000001001_0000000000000000;
      patterns[167] = 50'b11_0000000000000010_0000000000001001_0000000000001011;
      patterns[168] = 50'b00_0000000000000010_0000000000001010_0000000000001100;
      patterns[169] = 50'b01_0000000000000010_0000000000001010_1111111111111000;
      patterns[170] = 50'b10_0000000000000010_0000000000001010_0000000000000010;
      patterns[171] = 50'b11_0000000000000010_0000000000001010_0000000000001010;
      patterns[172] = 50'b00_0000000000000010_0000000000001011_0000000000001101;
      patterns[173] = 50'b01_0000000000000010_0000000000001011_1111111111110111;
      patterns[174] = 50'b10_0000000000000010_0000000000001011_0000000000000010;
      patterns[175] = 50'b11_0000000000000010_0000000000001011_0000000000001011;
      patterns[176] = 50'b00_0000000000000010_0000000000001100_0000000000001110;
      patterns[177] = 50'b01_0000000000000010_0000000000001100_1111111111110110;
      patterns[178] = 50'b10_0000000000000010_0000000000001100_0000000000000000;
      patterns[179] = 50'b11_0000000000000010_0000000000001100_0000000000001110;
      patterns[180] = 50'b00_0000000000000010_0000000000001101_0000000000001111;
      patterns[181] = 50'b01_0000000000000010_0000000000001101_1111111111110101;
      patterns[182] = 50'b10_0000000000000010_0000000000001101_0000000000000000;
      patterns[183] = 50'b11_0000000000000010_0000000000001101_0000000000001111;
      patterns[184] = 50'b00_0000000000000010_0000000000001110_0000000000010000;
      patterns[185] = 50'b01_0000000000000010_0000000000001110_1111111111110100;
      patterns[186] = 50'b10_0000000000000010_0000000000001110_0000000000000010;
      patterns[187] = 50'b11_0000000000000010_0000000000001110_0000000000001110;
      patterns[188] = 50'b00_0000000000000010_0000000000001111_0000000000010001;
      patterns[189] = 50'b01_0000000000000010_0000000000001111_1111111111110011;
      patterns[190] = 50'b10_0000000000000010_0000000000001111_0000000000000010;
      patterns[191] = 50'b11_0000000000000010_0000000000001111_0000000000001111;
      patterns[192] = 50'b00_0000000000000011_0000000000000000_0000000000000011;
      patterns[193] = 50'b01_0000000000000011_0000000000000000_0000000000000011;
      patterns[194] = 50'b10_0000000000000011_0000000000000000_0000000000000000;
      patterns[195] = 50'b11_0000000000000011_0000000000000000_0000000000000011;
      patterns[196] = 50'b00_0000000000000011_0000000000000001_0000000000000100;
      patterns[197] = 50'b01_0000000000000011_0000000000000001_0000000000000010;
      patterns[198] = 50'b10_0000000000000011_0000000000000001_0000000000000001;
      patterns[199] = 50'b11_0000000000000011_0000000000000001_0000000000000011;
      patterns[200] = 50'b00_0000000000000011_0000000000000010_0000000000000101;
      patterns[201] = 50'b01_0000000000000011_0000000000000010_0000000000000001;
      patterns[202] = 50'b10_0000000000000011_0000000000000010_0000000000000010;
      patterns[203] = 50'b11_0000000000000011_0000000000000010_0000000000000011;
      patterns[204] = 50'b00_0000000000000011_0000000000000011_0000000000000110;
      patterns[205] = 50'b01_0000000000000011_0000000000000011_0000000000000000;
      patterns[206] = 50'b10_0000000000000011_0000000000000011_0000000000000011;
      patterns[207] = 50'b11_0000000000000011_0000000000000011_0000000000000011;
      patterns[208] = 50'b00_0000000000000011_0000000000000100_0000000000000111;
      patterns[209] = 50'b01_0000000000000011_0000000000000100_1111111111111111;
      patterns[210] = 50'b10_0000000000000011_0000000000000100_0000000000000000;
      patterns[211] = 50'b11_0000000000000011_0000000000000100_0000000000000111;
      patterns[212] = 50'b00_0000000000000011_0000000000000101_0000000000001000;
      patterns[213] = 50'b01_0000000000000011_0000000000000101_1111111111111110;
      patterns[214] = 50'b10_0000000000000011_0000000000000101_0000000000000001;
      patterns[215] = 50'b11_0000000000000011_0000000000000101_0000000000000111;
      patterns[216] = 50'b00_0000000000000011_0000000000000110_0000000000001001;
      patterns[217] = 50'b01_0000000000000011_0000000000000110_1111111111111101;
      patterns[218] = 50'b10_0000000000000011_0000000000000110_0000000000000010;
      patterns[219] = 50'b11_0000000000000011_0000000000000110_0000000000000111;
      patterns[220] = 50'b00_0000000000000011_0000000000000111_0000000000001010;
      patterns[221] = 50'b01_0000000000000011_0000000000000111_1111111111111100;
      patterns[222] = 50'b10_0000000000000011_0000000000000111_0000000000000011;
      patterns[223] = 50'b11_0000000000000011_0000000000000111_0000000000000111;
      patterns[224] = 50'b00_0000000000000011_0000000000001000_0000000000001011;
      patterns[225] = 50'b01_0000000000000011_0000000000001000_1111111111111011;
      patterns[226] = 50'b10_0000000000000011_0000000000001000_0000000000000000;
      patterns[227] = 50'b11_0000000000000011_0000000000001000_0000000000001011;
      patterns[228] = 50'b00_0000000000000011_0000000000001001_0000000000001100;
      patterns[229] = 50'b01_0000000000000011_0000000000001001_1111111111111010;
      patterns[230] = 50'b10_0000000000000011_0000000000001001_0000000000000001;
      patterns[231] = 50'b11_0000000000000011_0000000000001001_0000000000001011;
      patterns[232] = 50'b00_0000000000000011_0000000000001010_0000000000001101;
      patterns[233] = 50'b01_0000000000000011_0000000000001010_1111111111111001;
      patterns[234] = 50'b10_0000000000000011_0000000000001010_0000000000000010;
      patterns[235] = 50'b11_0000000000000011_0000000000001010_0000000000001011;
      patterns[236] = 50'b00_0000000000000011_0000000000001011_0000000000001110;
      patterns[237] = 50'b01_0000000000000011_0000000000001011_1111111111111000;
      patterns[238] = 50'b10_0000000000000011_0000000000001011_0000000000000011;
      patterns[239] = 50'b11_0000000000000011_0000000000001011_0000000000001011;
      patterns[240] = 50'b00_0000000000000011_0000000000001100_0000000000001111;
      patterns[241] = 50'b01_0000000000000011_0000000000001100_1111111111110111;
      patterns[242] = 50'b10_0000000000000011_0000000000001100_0000000000000000;
      patterns[243] = 50'b11_0000000000000011_0000000000001100_0000000000001111;
      patterns[244] = 50'b00_0000000000000011_0000000000001101_0000000000010000;
      patterns[245] = 50'b01_0000000000000011_0000000000001101_1111111111110110;
      patterns[246] = 50'b10_0000000000000011_0000000000001101_0000000000000001;
      patterns[247] = 50'b11_0000000000000011_0000000000001101_0000000000001111;
      patterns[248] = 50'b00_0000000000000011_0000000000001110_0000000000010001;
      patterns[249] = 50'b01_0000000000000011_0000000000001110_1111111111110101;
      patterns[250] = 50'b10_0000000000000011_0000000000001110_0000000000000010;
      patterns[251] = 50'b11_0000000000000011_0000000000001110_0000000000001111;
      patterns[252] = 50'b00_0000000000000011_0000000000001111_0000000000010010;
      patterns[253] = 50'b01_0000000000000011_0000000000001111_1111111111110100;
      patterns[254] = 50'b10_0000000000000011_0000000000001111_0000000000000011;
      patterns[255] = 50'b11_0000000000000011_0000000000001111_0000000000001111;
      patterns[256] = 50'b00_0000000000000100_0000000000000000_0000000000000100;
      patterns[257] = 50'b01_0000000000000100_0000000000000000_0000000000000100;
      patterns[258] = 50'b10_0000000000000100_0000000000000000_0000000000000000;
      patterns[259] = 50'b11_0000000000000100_0000000000000000_0000000000000100;
      patterns[260] = 50'b00_0000000000000100_0000000000000001_0000000000000101;
      patterns[261] = 50'b01_0000000000000100_0000000000000001_0000000000000011;
      patterns[262] = 50'b10_0000000000000100_0000000000000001_0000000000000000;
      patterns[263] = 50'b11_0000000000000100_0000000000000001_0000000000000101;
      patterns[264] = 50'b00_0000000000000100_0000000000000010_0000000000000110;
      patterns[265] = 50'b01_0000000000000100_0000000000000010_0000000000000010;
      patterns[266] = 50'b10_0000000000000100_0000000000000010_0000000000000000;
      patterns[267] = 50'b11_0000000000000100_0000000000000010_0000000000000110;
      patterns[268] = 50'b00_0000000000000100_0000000000000011_0000000000000111;
      patterns[269] = 50'b01_0000000000000100_0000000000000011_0000000000000001;
      patterns[270] = 50'b10_0000000000000100_0000000000000011_0000000000000000;
      patterns[271] = 50'b11_0000000000000100_0000000000000011_0000000000000111;
      patterns[272] = 50'b00_0000000000000100_0000000000000100_0000000000001000;
      patterns[273] = 50'b01_0000000000000100_0000000000000100_0000000000000000;
      patterns[274] = 50'b10_0000000000000100_0000000000000100_0000000000000100;
      patterns[275] = 50'b11_0000000000000100_0000000000000100_0000000000000100;
      patterns[276] = 50'b00_0000000000000100_0000000000000101_0000000000001001;
      patterns[277] = 50'b01_0000000000000100_0000000000000101_1111111111111111;
      patterns[278] = 50'b10_0000000000000100_0000000000000101_0000000000000100;
      patterns[279] = 50'b11_0000000000000100_0000000000000101_0000000000000101;
      patterns[280] = 50'b00_0000000000000100_0000000000000110_0000000000001010;
      patterns[281] = 50'b01_0000000000000100_0000000000000110_1111111111111110;
      patterns[282] = 50'b10_0000000000000100_0000000000000110_0000000000000100;
      patterns[283] = 50'b11_0000000000000100_0000000000000110_0000000000000110;
      patterns[284] = 50'b00_0000000000000100_0000000000000111_0000000000001011;
      patterns[285] = 50'b01_0000000000000100_0000000000000111_1111111111111101;
      patterns[286] = 50'b10_0000000000000100_0000000000000111_0000000000000100;
      patterns[287] = 50'b11_0000000000000100_0000000000000111_0000000000000111;
      patterns[288] = 50'b00_0000000000000100_0000000000001000_0000000000001100;
      patterns[289] = 50'b01_0000000000000100_0000000000001000_1111111111111100;
      patterns[290] = 50'b10_0000000000000100_0000000000001000_0000000000000000;
      patterns[291] = 50'b11_0000000000000100_0000000000001000_0000000000001100;
      patterns[292] = 50'b00_0000000000000100_0000000000001001_0000000000001101;
      patterns[293] = 50'b01_0000000000000100_0000000000001001_1111111111111011;
      patterns[294] = 50'b10_0000000000000100_0000000000001001_0000000000000000;
      patterns[295] = 50'b11_0000000000000100_0000000000001001_0000000000001101;
      patterns[296] = 50'b00_0000000000000100_0000000000001010_0000000000001110;
      patterns[297] = 50'b01_0000000000000100_0000000000001010_1111111111111010;
      patterns[298] = 50'b10_0000000000000100_0000000000001010_0000000000000000;
      patterns[299] = 50'b11_0000000000000100_0000000000001010_0000000000001110;
      patterns[300] = 50'b00_0000000000000100_0000000000001011_0000000000001111;
      patterns[301] = 50'b01_0000000000000100_0000000000001011_1111111111111001;
      patterns[302] = 50'b10_0000000000000100_0000000000001011_0000000000000000;
      patterns[303] = 50'b11_0000000000000100_0000000000001011_0000000000001111;
      patterns[304] = 50'b00_0000000000000100_0000000000001100_0000000000010000;
      patterns[305] = 50'b01_0000000000000100_0000000000001100_1111111111111000;
      patterns[306] = 50'b10_0000000000000100_0000000000001100_0000000000000100;
      patterns[307] = 50'b11_0000000000000100_0000000000001100_0000000000001100;
      patterns[308] = 50'b00_0000000000000100_0000000000001101_0000000000010001;
      patterns[309] = 50'b01_0000000000000100_0000000000001101_1111111111110111;
      patterns[310] = 50'b10_0000000000000100_0000000000001101_0000000000000100;
      patterns[311] = 50'b11_0000000000000100_0000000000001101_0000000000001101;
      patterns[312] = 50'b00_0000000000000100_0000000000001110_0000000000010010;
      patterns[313] = 50'b01_0000000000000100_0000000000001110_1111111111110110;
      patterns[314] = 50'b10_0000000000000100_0000000000001110_0000000000000100;
      patterns[315] = 50'b11_0000000000000100_0000000000001110_0000000000001110;
      patterns[316] = 50'b00_0000000000000100_0000000000001111_0000000000010011;
      patterns[317] = 50'b01_0000000000000100_0000000000001111_1111111111110101;
      patterns[318] = 50'b10_0000000000000100_0000000000001111_0000000000000100;
      patterns[319] = 50'b11_0000000000000100_0000000000001111_0000000000001111;
      patterns[320] = 50'b00_0000000000000101_0000000000000000_0000000000000101;
      patterns[321] = 50'b01_0000000000000101_0000000000000000_0000000000000101;
      patterns[322] = 50'b10_0000000000000101_0000000000000000_0000000000000000;
      patterns[323] = 50'b11_0000000000000101_0000000000000000_0000000000000101;
      patterns[324] = 50'b00_0000000000000101_0000000000000001_0000000000000110;
      patterns[325] = 50'b01_0000000000000101_0000000000000001_0000000000000100;
      patterns[326] = 50'b10_0000000000000101_0000000000000001_0000000000000001;
      patterns[327] = 50'b11_0000000000000101_0000000000000001_0000000000000101;
      patterns[328] = 50'b00_0000000000000101_0000000000000010_0000000000000111;
      patterns[329] = 50'b01_0000000000000101_0000000000000010_0000000000000011;
      patterns[330] = 50'b10_0000000000000101_0000000000000010_0000000000000000;
      patterns[331] = 50'b11_0000000000000101_0000000000000010_0000000000000111;
      patterns[332] = 50'b00_0000000000000101_0000000000000011_0000000000001000;
      patterns[333] = 50'b01_0000000000000101_0000000000000011_0000000000000010;
      patterns[334] = 50'b10_0000000000000101_0000000000000011_0000000000000001;
      patterns[335] = 50'b11_0000000000000101_0000000000000011_0000000000000111;
      patterns[336] = 50'b00_0000000000000101_0000000000000100_0000000000001001;
      patterns[337] = 50'b01_0000000000000101_0000000000000100_0000000000000001;
      patterns[338] = 50'b10_0000000000000101_0000000000000100_0000000000000100;
      patterns[339] = 50'b11_0000000000000101_0000000000000100_0000000000000101;
      patterns[340] = 50'b00_0000000000000101_0000000000000101_0000000000001010;
      patterns[341] = 50'b01_0000000000000101_0000000000000101_0000000000000000;
      patterns[342] = 50'b10_0000000000000101_0000000000000101_0000000000000101;
      patterns[343] = 50'b11_0000000000000101_0000000000000101_0000000000000101;
      patterns[344] = 50'b00_0000000000000101_0000000000000110_0000000000001011;
      patterns[345] = 50'b01_0000000000000101_0000000000000110_1111111111111111;
      patterns[346] = 50'b10_0000000000000101_0000000000000110_0000000000000100;
      patterns[347] = 50'b11_0000000000000101_0000000000000110_0000000000000111;
      patterns[348] = 50'b00_0000000000000101_0000000000000111_0000000000001100;
      patterns[349] = 50'b01_0000000000000101_0000000000000111_1111111111111110;
      patterns[350] = 50'b10_0000000000000101_0000000000000111_0000000000000101;
      patterns[351] = 50'b11_0000000000000101_0000000000000111_0000000000000111;
      patterns[352] = 50'b00_0000000000000101_0000000000001000_0000000000001101;
      patterns[353] = 50'b01_0000000000000101_0000000000001000_1111111111111101;
      patterns[354] = 50'b10_0000000000000101_0000000000001000_0000000000000000;
      patterns[355] = 50'b11_0000000000000101_0000000000001000_0000000000001101;
      patterns[356] = 50'b00_0000000000000101_0000000000001001_0000000000001110;
      patterns[357] = 50'b01_0000000000000101_0000000000001001_1111111111111100;
      patterns[358] = 50'b10_0000000000000101_0000000000001001_0000000000000001;
      patterns[359] = 50'b11_0000000000000101_0000000000001001_0000000000001101;
      patterns[360] = 50'b00_0000000000000101_0000000000001010_0000000000001111;
      patterns[361] = 50'b01_0000000000000101_0000000000001010_1111111111111011;
      patterns[362] = 50'b10_0000000000000101_0000000000001010_0000000000000000;
      patterns[363] = 50'b11_0000000000000101_0000000000001010_0000000000001111;
      patterns[364] = 50'b00_0000000000000101_0000000000001011_0000000000010000;
      patterns[365] = 50'b01_0000000000000101_0000000000001011_1111111111111010;
      patterns[366] = 50'b10_0000000000000101_0000000000001011_0000000000000001;
      patterns[367] = 50'b11_0000000000000101_0000000000001011_0000000000001111;
      patterns[368] = 50'b00_0000000000000101_0000000000001100_0000000000010001;
      patterns[369] = 50'b01_0000000000000101_0000000000001100_1111111111111001;
      patterns[370] = 50'b10_0000000000000101_0000000000001100_0000000000000100;
      patterns[371] = 50'b11_0000000000000101_0000000000001100_0000000000001101;
      patterns[372] = 50'b00_0000000000000101_0000000000001101_0000000000010010;
      patterns[373] = 50'b01_0000000000000101_0000000000001101_1111111111111000;
      patterns[374] = 50'b10_0000000000000101_0000000000001101_0000000000000101;
      patterns[375] = 50'b11_0000000000000101_0000000000001101_0000000000001101;
      patterns[376] = 50'b00_0000000000000101_0000000000001110_0000000000010011;
      patterns[377] = 50'b01_0000000000000101_0000000000001110_1111111111110111;
      patterns[378] = 50'b10_0000000000000101_0000000000001110_0000000000000100;
      patterns[379] = 50'b11_0000000000000101_0000000000001110_0000000000001111;
      patterns[380] = 50'b00_0000000000000101_0000000000001111_0000000000010100;
      patterns[381] = 50'b01_0000000000000101_0000000000001111_1111111111110110;
      patterns[382] = 50'b10_0000000000000101_0000000000001111_0000000000000101;
      patterns[383] = 50'b11_0000000000000101_0000000000001111_0000000000001111;
      patterns[384] = 50'b00_0000000000000110_0000000000000000_0000000000000110;
      patterns[385] = 50'b01_0000000000000110_0000000000000000_0000000000000110;
      patterns[386] = 50'b10_0000000000000110_0000000000000000_0000000000000000;
      patterns[387] = 50'b11_0000000000000110_0000000000000000_0000000000000110;
      patterns[388] = 50'b00_0000000000000110_0000000000000001_0000000000000111;
      patterns[389] = 50'b01_0000000000000110_0000000000000001_0000000000000101;
      patterns[390] = 50'b10_0000000000000110_0000000000000001_0000000000000000;
      patterns[391] = 50'b11_0000000000000110_0000000000000001_0000000000000111;
      patterns[392] = 50'b00_0000000000000110_0000000000000010_0000000000001000;
      patterns[393] = 50'b01_0000000000000110_0000000000000010_0000000000000100;
      patterns[394] = 50'b10_0000000000000110_0000000000000010_0000000000000010;
      patterns[395] = 50'b11_0000000000000110_0000000000000010_0000000000000110;
      patterns[396] = 50'b00_0000000000000110_0000000000000011_0000000000001001;
      patterns[397] = 50'b01_0000000000000110_0000000000000011_0000000000000011;
      patterns[398] = 50'b10_0000000000000110_0000000000000011_0000000000000010;
      patterns[399] = 50'b11_0000000000000110_0000000000000011_0000000000000111;
      patterns[400] = 50'b00_0000000000000110_0000000000000100_0000000000001010;
      patterns[401] = 50'b01_0000000000000110_0000000000000100_0000000000000010;
      patterns[402] = 50'b10_0000000000000110_0000000000000100_0000000000000100;
      patterns[403] = 50'b11_0000000000000110_0000000000000100_0000000000000110;
      patterns[404] = 50'b00_0000000000000110_0000000000000101_0000000000001011;
      patterns[405] = 50'b01_0000000000000110_0000000000000101_0000000000000001;
      patterns[406] = 50'b10_0000000000000110_0000000000000101_0000000000000100;
      patterns[407] = 50'b11_0000000000000110_0000000000000101_0000000000000111;
      patterns[408] = 50'b00_0000000000000110_0000000000000110_0000000000001100;
      patterns[409] = 50'b01_0000000000000110_0000000000000110_0000000000000000;
      patterns[410] = 50'b10_0000000000000110_0000000000000110_0000000000000110;
      patterns[411] = 50'b11_0000000000000110_0000000000000110_0000000000000110;
      patterns[412] = 50'b00_0000000000000110_0000000000000111_0000000000001101;
      patterns[413] = 50'b01_0000000000000110_0000000000000111_1111111111111111;
      patterns[414] = 50'b10_0000000000000110_0000000000000111_0000000000000110;
      patterns[415] = 50'b11_0000000000000110_0000000000000111_0000000000000111;
      patterns[416] = 50'b00_0000000000000110_0000000000001000_0000000000001110;
      patterns[417] = 50'b01_0000000000000110_0000000000001000_1111111111111110;
      patterns[418] = 50'b10_0000000000000110_0000000000001000_0000000000000000;
      patterns[419] = 50'b11_0000000000000110_0000000000001000_0000000000001110;
      patterns[420] = 50'b00_0000000000000110_0000000000001001_0000000000001111;
      patterns[421] = 50'b01_0000000000000110_0000000000001001_1111111111111101;
      patterns[422] = 50'b10_0000000000000110_0000000000001001_0000000000000000;
      patterns[423] = 50'b11_0000000000000110_0000000000001001_0000000000001111;
      patterns[424] = 50'b00_0000000000000110_0000000000001010_0000000000010000;
      patterns[425] = 50'b01_0000000000000110_0000000000001010_1111111111111100;
      patterns[426] = 50'b10_0000000000000110_0000000000001010_0000000000000010;
      patterns[427] = 50'b11_0000000000000110_0000000000001010_0000000000001110;
      patterns[428] = 50'b00_0000000000000110_0000000000001011_0000000000010001;
      patterns[429] = 50'b01_0000000000000110_0000000000001011_1111111111111011;
      patterns[430] = 50'b10_0000000000000110_0000000000001011_0000000000000010;
      patterns[431] = 50'b11_0000000000000110_0000000000001011_0000000000001111;
      patterns[432] = 50'b00_0000000000000110_0000000000001100_0000000000010010;
      patterns[433] = 50'b01_0000000000000110_0000000000001100_1111111111111010;
      patterns[434] = 50'b10_0000000000000110_0000000000001100_0000000000000100;
      patterns[435] = 50'b11_0000000000000110_0000000000001100_0000000000001110;
      patterns[436] = 50'b00_0000000000000110_0000000000001101_0000000000010011;
      patterns[437] = 50'b01_0000000000000110_0000000000001101_1111111111111001;
      patterns[438] = 50'b10_0000000000000110_0000000000001101_0000000000000100;
      patterns[439] = 50'b11_0000000000000110_0000000000001101_0000000000001111;
      patterns[440] = 50'b00_0000000000000110_0000000000001110_0000000000010100;
      patterns[441] = 50'b01_0000000000000110_0000000000001110_1111111111111000;
      patterns[442] = 50'b10_0000000000000110_0000000000001110_0000000000000110;
      patterns[443] = 50'b11_0000000000000110_0000000000001110_0000000000001110;
      patterns[444] = 50'b00_0000000000000110_0000000000001111_0000000000010101;
      patterns[445] = 50'b01_0000000000000110_0000000000001111_1111111111110111;
      patterns[446] = 50'b10_0000000000000110_0000000000001111_0000000000000110;
      patterns[447] = 50'b11_0000000000000110_0000000000001111_0000000000001111;
      patterns[448] = 50'b00_0000000000000111_0000000000000000_0000000000000111;
      patterns[449] = 50'b01_0000000000000111_0000000000000000_0000000000000111;
      patterns[450] = 50'b10_0000000000000111_0000000000000000_0000000000000000;
      patterns[451] = 50'b11_0000000000000111_0000000000000000_0000000000000111;
      patterns[452] = 50'b00_0000000000000111_0000000000000001_0000000000001000;
      patterns[453] = 50'b01_0000000000000111_0000000000000001_0000000000000110;
      patterns[454] = 50'b10_0000000000000111_0000000000000001_0000000000000001;
      patterns[455] = 50'b11_0000000000000111_0000000000000001_0000000000000111;
      patterns[456] = 50'b00_0000000000000111_0000000000000010_0000000000001001;
      patterns[457] = 50'b01_0000000000000111_0000000000000010_0000000000000101;
      patterns[458] = 50'b10_0000000000000111_0000000000000010_0000000000000010;
      patterns[459] = 50'b11_0000000000000111_0000000000000010_0000000000000111;
      patterns[460] = 50'b00_0000000000000111_0000000000000011_0000000000001010;
      patterns[461] = 50'b01_0000000000000111_0000000000000011_0000000000000100;
      patterns[462] = 50'b10_0000000000000111_0000000000000011_0000000000000011;
      patterns[463] = 50'b11_0000000000000111_0000000000000011_0000000000000111;
      patterns[464] = 50'b00_0000000000000111_0000000000000100_0000000000001011;
      patterns[465] = 50'b01_0000000000000111_0000000000000100_0000000000000011;
      patterns[466] = 50'b10_0000000000000111_0000000000000100_0000000000000100;
      patterns[467] = 50'b11_0000000000000111_0000000000000100_0000000000000111;
      patterns[468] = 50'b00_0000000000000111_0000000000000101_0000000000001100;
      patterns[469] = 50'b01_0000000000000111_0000000000000101_0000000000000010;
      patterns[470] = 50'b10_0000000000000111_0000000000000101_0000000000000101;
      patterns[471] = 50'b11_0000000000000111_0000000000000101_0000000000000111;
      patterns[472] = 50'b00_0000000000000111_0000000000000110_0000000000001101;
      patterns[473] = 50'b01_0000000000000111_0000000000000110_0000000000000001;
      patterns[474] = 50'b10_0000000000000111_0000000000000110_0000000000000110;
      patterns[475] = 50'b11_0000000000000111_0000000000000110_0000000000000111;
      patterns[476] = 50'b00_0000000000000111_0000000000000111_0000000000001110;
      patterns[477] = 50'b01_0000000000000111_0000000000000111_0000000000000000;
      patterns[478] = 50'b10_0000000000000111_0000000000000111_0000000000000111;
      patterns[479] = 50'b11_0000000000000111_0000000000000111_0000000000000111;
      patterns[480] = 50'b00_0000000000000111_0000000000001000_0000000000001111;
      patterns[481] = 50'b01_0000000000000111_0000000000001000_1111111111111111;
      patterns[482] = 50'b10_0000000000000111_0000000000001000_0000000000000000;
      patterns[483] = 50'b11_0000000000000111_0000000000001000_0000000000001111;
      patterns[484] = 50'b00_0000000000000111_0000000000001001_0000000000010000;
      patterns[485] = 50'b01_0000000000000111_0000000000001001_1111111111111110;
      patterns[486] = 50'b10_0000000000000111_0000000000001001_0000000000000001;
      patterns[487] = 50'b11_0000000000000111_0000000000001001_0000000000001111;
      patterns[488] = 50'b00_0000000000000111_0000000000001010_0000000000010001;
      patterns[489] = 50'b01_0000000000000111_0000000000001010_1111111111111101;
      patterns[490] = 50'b10_0000000000000111_0000000000001010_0000000000000010;
      patterns[491] = 50'b11_0000000000000111_0000000000001010_0000000000001111;
      patterns[492] = 50'b00_0000000000000111_0000000000001011_0000000000010010;
      patterns[493] = 50'b01_0000000000000111_0000000000001011_1111111111111100;
      patterns[494] = 50'b10_0000000000000111_0000000000001011_0000000000000011;
      patterns[495] = 50'b11_0000000000000111_0000000000001011_0000000000001111;
      patterns[496] = 50'b00_0000000000000111_0000000000001100_0000000000010011;
      patterns[497] = 50'b01_0000000000000111_0000000000001100_1111111111111011;
      patterns[498] = 50'b10_0000000000000111_0000000000001100_0000000000000100;
      patterns[499] = 50'b11_0000000000000111_0000000000001100_0000000000001111;
      patterns[500] = 50'b00_0000000000000111_0000000000001101_0000000000010100;
      patterns[501] = 50'b01_0000000000000111_0000000000001101_1111111111111010;
      patterns[502] = 50'b10_0000000000000111_0000000000001101_0000000000000101;
      patterns[503] = 50'b11_0000000000000111_0000000000001101_0000000000001111;
      patterns[504] = 50'b00_0000000000000111_0000000000001110_0000000000010101;
      patterns[505] = 50'b01_0000000000000111_0000000000001110_1111111111111001;
      patterns[506] = 50'b10_0000000000000111_0000000000001110_0000000000000110;
      patterns[507] = 50'b11_0000000000000111_0000000000001110_0000000000001111;
      patterns[508] = 50'b00_0000000000000111_0000000000001111_0000000000010110;
      patterns[509] = 50'b01_0000000000000111_0000000000001111_1111111111111000;
      patterns[510] = 50'b10_0000000000000111_0000000000001111_0000000000000111;
      patterns[511] = 50'b11_0000000000000111_0000000000001111_0000000000001111;
      patterns[512] = 50'b00_0000000000001000_0000000000000000_0000000000001000;
      patterns[513] = 50'b01_0000000000001000_0000000000000000_0000000000001000;
      patterns[514] = 50'b10_0000000000001000_0000000000000000_0000000000000000;
      patterns[515] = 50'b11_0000000000001000_0000000000000000_0000000000001000;
      patterns[516] = 50'b00_0000000000001000_0000000000000001_0000000000001001;
      patterns[517] = 50'b01_0000000000001000_0000000000000001_0000000000000111;
      patterns[518] = 50'b10_0000000000001000_0000000000000001_0000000000000000;
      patterns[519] = 50'b11_0000000000001000_0000000000000001_0000000000001001;
      patterns[520] = 50'b00_0000000000001000_0000000000000010_0000000000001010;
      patterns[521] = 50'b01_0000000000001000_0000000000000010_0000000000000110;
      patterns[522] = 50'b10_0000000000001000_0000000000000010_0000000000000000;
      patterns[523] = 50'b11_0000000000001000_0000000000000010_0000000000001010;
      patterns[524] = 50'b00_0000000000001000_0000000000000011_0000000000001011;
      patterns[525] = 50'b01_0000000000001000_0000000000000011_0000000000000101;
      patterns[526] = 50'b10_0000000000001000_0000000000000011_0000000000000000;
      patterns[527] = 50'b11_0000000000001000_0000000000000011_0000000000001011;
      patterns[528] = 50'b00_0000000000001000_0000000000000100_0000000000001100;
      patterns[529] = 50'b01_0000000000001000_0000000000000100_0000000000000100;
      patterns[530] = 50'b10_0000000000001000_0000000000000100_0000000000000000;
      patterns[531] = 50'b11_0000000000001000_0000000000000100_0000000000001100;
      patterns[532] = 50'b00_0000000000001000_0000000000000101_0000000000001101;
      patterns[533] = 50'b01_0000000000001000_0000000000000101_0000000000000011;
      patterns[534] = 50'b10_0000000000001000_0000000000000101_0000000000000000;
      patterns[535] = 50'b11_0000000000001000_0000000000000101_0000000000001101;
      patterns[536] = 50'b00_0000000000001000_0000000000000110_0000000000001110;
      patterns[537] = 50'b01_0000000000001000_0000000000000110_0000000000000010;
      patterns[538] = 50'b10_0000000000001000_0000000000000110_0000000000000000;
      patterns[539] = 50'b11_0000000000001000_0000000000000110_0000000000001110;
      patterns[540] = 50'b00_0000000000001000_0000000000000111_0000000000001111;
      patterns[541] = 50'b01_0000000000001000_0000000000000111_0000000000000001;
      patterns[542] = 50'b10_0000000000001000_0000000000000111_0000000000000000;
      patterns[543] = 50'b11_0000000000001000_0000000000000111_0000000000001111;
      patterns[544] = 50'b00_0000000000001000_0000000000001000_0000000000010000;
      patterns[545] = 50'b01_0000000000001000_0000000000001000_0000000000000000;
      patterns[546] = 50'b10_0000000000001000_0000000000001000_0000000000001000;
      patterns[547] = 50'b11_0000000000001000_0000000000001000_0000000000001000;
      patterns[548] = 50'b00_0000000000001000_0000000000001001_0000000000010001;
      patterns[549] = 50'b01_0000000000001000_0000000000001001_1111111111111111;
      patterns[550] = 50'b10_0000000000001000_0000000000001001_0000000000001000;
      patterns[551] = 50'b11_0000000000001000_0000000000001001_0000000000001001;
      patterns[552] = 50'b00_0000000000001000_0000000000001010_0000000000010010;
      patterns[553] = 50'b01_0000000000001000_0000000000001010_1111111111111110;
      patterns[554] = 50'b10_0000000000001000_0000000000001010_0000000000001000;
      patterns[555] = 50'b11_0000000000001000_0000000000001010_0000000000001010;
      patterns[556] = 50'b00_0000000000001000_0000000000001011_0000000000010011;
      patterns[557] = 50'b01_0000000000001000_0000000000001011_1111111111111101;
      patterns[558] = 50'b10_0000000000001000_0000000000001011_0000000000001000;
      patterns[559] = 50'b11_0000000000001000_0000000000001011_0000000000001011;
      patterns[560] = 50'b00_0000000000001000_0000000000001100_0000000000010100;
      patterns[561] = 50'b01_0000000000001000_0000000000001100_1111111111111100;
      patterns[562] = 50'b10_0000000000001000_0000000000001100_0000000000001000;
      patterns[563] = 50'b11_0000000000001000_0000000000001100_0000000000001100;
      patterns[564] = 50'b00_0000000000001000_0000000000001101_0000000000010101;
      patterns[565] = 50'b01_0000000000001000_0000000000001101_1111111111111011;
      patterns[566] = 50'b10_0000000000001000_0000000000001101_0000000000001000;
      patterns[567] = 50'b11_0000000000001000_0000000000001101_0000000000001101;
      patterns[568] = 50'b00_0000000000001000_0000000000001110_0000000000010110;
      patterns[569] = 50'b01_0000000000001000_0000000000001110_1111111111111010;
      patterns[570] = 50'b10_0000000000001000_0000000000001110_0000000000001000;
      patterns[571] = 50'b11_0000000000001000_0000000000001110_0000000000001110;
      patterns[572] = 50'b00_0000000000001000_0000000000001111_0000000000010111;
      patterns[573] = 50'b01_0000000000001000_0000000000001111_1111111111111001;
      patterns[574] = 50'b10_0000000000001000_0000000000001111_0000000000001000;
      patterns[575] = 50'b11_0000000000001000_0000000000001111_0000000000001111;
      patterns[576] = 50'b00_0000000000001001_0000000000000000_0000000000001001;
      patterns[577] = 50'b01_0000000000001001_0000000000000000_0000000000001001;
      patterns[578] = 50'b10_0000000000001001_0000000000000000_0000000000000000;
      patterns[579] = 50'b11_0000000000001001_0000000000000000_0000000000001001;
      patterns[580] = 50'b00_0000000000001001_0000000000000001_0000000000001010;
      patterns[581] = 50'b01_0000000000001001_0000000000000001_0000000000001000;
      patterns[582] = 50'b10_0000000000001001_0000000000000001_0000000000000001;
      patterns[583] = 50'b11_0000000000001001_0000000000000001_0000000000001001;
      patterns[584] = 50'b00_0000000000001001_0000000000000010_0000000000001011;
      patterns[585] = 50'b01_0000000000001001_0000000000000010_0000000000000111;
      patterns[586] = 50'b10_0000000000001001_0000000000000010_0000000000000000;
      patterns[587] = 50'b11_0000000000001001_0000000000000010_0000000000001011;
      patterns[588] = 50'b00_0000000000001001_0000000000000011_0000000000001100;
      patterns[589] = 50'b01_0000000000001001_0000000000000011_0000000000000110;
      patterns[590] = 50'b10_0000000000001001_0000000000000011_0000000000000001;
      patterns[591] = 50'b11_0000000000001001_0000000000000011_0000000000001011;
      patterns[592] = 50'b00_0000000000001001_0000000000000100_0000000000001101;
      patterns[593] = 50'b01_0000000000001001_0000000000000100_0000000000000101;
      patterns[594] = 50'b10_0000000000001001_0000000000000100_0000000000000000;
      patterns[595] = 50'b11_0000000000001001_0000000000000100_0000000000001101;
      patterns[596] = 50'b00_0000000000001001_0000000000000101_0000000000001110;
      patterns[597] = 50'b01_0000000000001001_0000000000000101_0000000000000100;
      patterns[598] = 50'b10_0000000000001001_0000000000000101_0000000000000001;
      patterns[599] = 50'b11_0000000000001001_0000000000000101_0000000000001101;
      patterns[600] = 50'b00_0000000000001001_0000000000000110_0000000000001111;
      patterns[601] = 50'b01_0000000000001001_0000000000000110_0000000000000011;
      patterns[602] = 50'b10_0000000000001001_0000000000000110_0000000000000000;
      patterns[603] = 50'b11_0000000000001001_0000000000000110_0000000000001111;
      patterns[604] = 50'b00_0000000000001001_0000000000000111_0000000000010000;
      patterns[605] = 50'b01_0000000000001001_0000000000000111_0000000000000010;
      patterns[606] = 50'b10_0000000000001001_0000000000000111_0000000000000001;
      patterns[607] = 50'b11_0000000000001001_0000000000000111_0000000000001111;
      patterns[608] = 50'b00_0000000000001001_0000000000001000_0000000000010001;
      patterns[609] = 50'b01_0000000000001001_0000000000001000_0000000000000001;
      patterns[610] = 50'b10_0000000000001001_0000000000001000_0000000000001000;
      patterns[611] = 50'b11_0000000000001001_0000000000001000_0000000000001001;
      patterns[612] = 50'b00_0000000000001001_0000000000001001_0000000000010010;
      patterns[613] = 50'b01_0000000000001001_0000000000001001_0000000000000000;
      patterns[614] = 50'b10_0000000000001001_0000000000001001_0000000000001001;
      patterns[615] = 50'b11_0000000000001001_0000000000001001_0000000000001001;
      patterns[616] = 50'b00_0000000000001001_0000000000001010_0000000000010011;
      patterns[617] = 50'b01_0000000000001001_0000000000001010_1111111111111111;
      patterns[618] = 50'b10_0000000000001001_0000000000001010_0000000000001000;
      patterns[619] = 50'b11_0000000000001001_0000000000001010_0000000000001011;
      patterns[620] = 50'b00_0000000000001001_0000000000001011_0000000000010100;
      patterns[621] = 50'b01_0000000000001001_0000000000001011_1111111111111110;
      patterns[622] = 50'b10_0000000000001001_0000000000001011_0000000000001001;
      patterns[623] = 50'b11_0000000000001001_0000000000001011_0000000000001011;
      patterns[624] = 50'b00_0000000000001001_0000000000001100_0000000000010101;
      patterns[625] = 50'b01_0000000000001001_0000000000001100_1111111111111101;
      patterns[626] = 50'b10_0000000000001001_0000000000001100_0000000000001000;
      patterns[627] = 50'b11_0000000000001001_0000000000001100_0000000000001101;
      patterns[628] = 50'b00_0000000000001001_0000000000001101_0000000000010110;
      patterns[629] = 50'b01_0000000000001001_0000000000001101_1111111111111100;
      patterns[630] = 50'b10_0000000000001001_0000000000001101_0000000000001001;
      patterns[631] = 50'b11_0000000000001001_0000000000001101_0000000000001101;
      patterns[632] = 50'b00_0000000000001001_0000000000001110_0000000000010111;
      patterns[633] = 50'b01_0000000000001001_0000000000001110_1111111111111011;
      patterns[634] = 50'b10_0000000000001001_0000000000001110_0000000000001000;
      patterns[635] = 50'b11_0000000000001001_0000000000001110_0000000000001111;
      patterns[636] = 50'b00_0000000000001001_0000000000001111_0000000000011000;
      patterns[637] = 50'b01_0000000000001001_0000000000001111_1111111111111010;
      patterns[638] = 50'b10_0000000000001001_0000000000001111_0000000000001001;
      patterns[639] = 50'b11_0000000000001001_0000000000001111_0000000000001111;
      patterns[640] = 50'b00_0000000000001010_0000000000000000_0000000000001010;
      patterns[641] = 50'b01_0000000000001010_0000000000000000_0000000000001010;
      patterns[642] = 50'b10_0000000000001010_0000000000000000_0000000000000000;
      patterns[643] = 50'b11_0000000000001010_0000000000000000_0000000000001010;
      patterns[644] = 50'b00_0000000000001010_0000000000000001_0000000000001011;
      patterns[645] = 50'b01_0000000000001010_0000000000000001_0000000000001001;
      patterns[646] = 50'b10_0000000000001010_0000000000000001_0000000000000000;
      patterns[647] = 50'b11_0000000000001010_0000000000000001_0000000000001011;
      patterns[648] = 50'b00_0000000000001010_0000000000000010_0000000000001100;
      patterns[649] = 50'b01_0000000000001010_0000000000000010_0000000000001000;
      patterns[650] = 50'b10_0000000000001010_0000000000000010_0000000000000010;
      patterns[651] = 50'b11_0000000000001010_0000000000000010_0000000000001010;
      patterns[652] = 50'b00_0000000000001010_0000000000000011_0000000000001101;
      patterns[653] = 50'b01_0000000000001010_0000000000000011_0000000000000111;
      patterns[654] = 50'b10_0000000000001010_0000000000000011_0000000000000010;
      patterns[655] = 50'b11_0000000000001010_0000000000000011_0000000000001011;
      patterns[656] = 50'b00_0000000000001010_0000000000000100_0000000000001110;
      patterns[657] = 50'b01_0000000000001010_0000000000000100_0000000000000110;
      patterns[658] = 50'b10_0000000000001010_0000000000000100_0000000000000000;
      patterns[659] = 50'b11_0000000000001010_0000000000000100_0000000000001110;
      patterns[660] = 50'b00_0000000000001010_0000000000000101_0000000000001111;
      patterns[661] = 50'b01_0000000000001010_0000000000000101_0000000000000101;
      patterns[662] = 50'b10_0000000000001010_0000000000000101_0000000000000000;
      patterns[663] = 50'b11_0000000000001010_0000000000000101_0000000000001111;
      patterns[664] = 50'b00_0000000000001010_0000000000000110_0000000000010000;
      patterns[665] = 50'b01_0000000000001010_0000000000000110_0000000000000100;
      patterns[666] = 50'b10_0000000000001010_0000000000000110_0000000000000010;
      patterns[667] = 50'b11_0000000000001010_0000000000000110_0000000000001110;
      patterns[668] = 50'b00_0000000000001010_0000000000000111_0000000000010001;
      patterns[669] = 50'b01_0000000000001010_0000000000000111_0000000000000011;
      patterns[670] = 50'b10_0000000000001010_0000000000000111_0000000000000010;
      patterns[671] = 50'b11_0000000000001010_0000000000000111_0000000000001111;
      patterns[672] = 50'b00_0000000000001010_0000000000001000_0000000000010010;
      patterns[673] = 50'b01_0000000000001010_0000000000001000_0000000000000010;
      patterns[674] = 50'b10_0000000000001010_0000000000001000_0000000000001000;
      patterns[675] = 50'b11_0000000000001010_0000000000001000_0000000000001010;
      patterns[676] = 50'b00_0000000000001010_0000000000001001_0000000000010011;
      patterns[677] = 50'b01_0000000000001010_0000000000001001_0000000000000001;
      patterns[678] = 50'b10_0000000000001010_0000000000001001_0000000000001000;
      patterns[679] = 50'b11_0000000000001010_0000000000001001_0000000000001011;
      patterns[680] = 50'b00_0000000000001010_0000000000001010_0000000000010100;
      patterns[681] = 50'b01_0000000000001010_0000000000001010_0000000000000000;
      patterns[682] = 50'b10_0000000000001010_0000000000001010_0000000000001010;
      patterns[683] = 50'b11_0000000000001010_0000000000001010_0000000000001010;
      patterns[684] = 50'b00_0000000000001010_0000000000001011_0000000000010101;
      patterns[685] = 50'b01_0000000000001010_0000000000001011_1111111111111111;
      patterns[686] = 50'b10_0000000000001010_0000000000001011_0000000000001010;
      patterns[687] = 50'b11_0000000000001010_0000000000001011_0000000000001011;
      patterns[688] = 50'b00_0000000000001010_0000000000001100_0000000000010110;
      patterns[689] = 50'b01_0000000000001010_0000000000001100_1111111111111110;
      patterns[690] = 50'b10_0000000000001010_0000000000001100_0000000000001000;
      patterns[691] = 50'b11_0000000000001010_0000000000001100_0000000000001110;
      patterns[692] = 50'b00_0000000000001010_0000000000001101_0000000000010111;
      patterns[693] = 50'b01_0000000000001010_0000000000001101_1111111111111101;
      patterns[694] = 50'b10_0000000000001010_0000000000001101_0000000000001000;
      patterns[695] = 50'b11_0000000000001010_0000000000001101_0000000000001111;
      patterns[696] = 50'b00_0000000000001010_0000000000001110_0000000000011000;
      patterns[697] = 50'b01_0000000000001010_0000000000001110_1111111111111100;
      patterns[698] = 50'b10_0000000000001010_0000000000001110_0000000000001010;
      patterns[699] = 50'b11_0000000000001010_0000000000001110_0000000000001110;
      patterns[700] = 50'b00_0000000000001010_0000000000001111_0000000000011001;
      patterns[701] = 50'b01_0000000000001010_0000000000001111_1111111111111011;
      patterns[702] = 50'b10_0000000000001010_0000000000001111_0000000000001010;
      patterns[703] = 50'b11_0000000000001010_0000000000001111_0000000000001111;
      patterns[704] = 50'b00_0000000000001011_0000000000000000_0000000000001011;
      patterns[705] = 50'b01_0000000000001011_0000000000000000_0000000000001011;
      patterns[706] = 50'b10_0000000000001011_0000000000000000_0000000000000000;
      patterns[707] = 50'b11_0000000000001011_0000000000000000_0000000000001011;
      patterns[708] = 50'b00_0000000000001011_0000000000000001_0000000000001100;
      patterns[709] = 50'b01_0000000000001011_0000000000000001_0000000000001010;
      patterns[710] = 50'b10_0000000000001011_0000000000000001_0000000000000001;
      patterns[711] = 50'b11_0000000000001011_0000000000000001_0000000000001011;
      patterns[712] = 50'b00_0000000000001011_0000000000000010_0000000000001101;
      patterns[713] = 50'b01_0000000000001011_0000000000000010_0000000000001001;
      patterns[714] = 50'b10_0000000000001011_0000000000000010_0000000000000010;
      patterns[715] = 50'b11_0000000000001011_0000000000000010_0000000000001011;
      patterns[716] = 50'b00_0000000000001011_0000000000000011_0000000000001110;
      patterns[717] = 50'b01_0000000000001011_0000000000000011_0000000000001000;
      patterns[718] = 50'b10_0000000000001011_0000000000000011_0000000000000011;
      patterns[719] = 50'b11_0000000000001011_0000000000000011_0000000000001011;
      patterns[720] = 50'b00_0000000000001011_0000000000000100_0000000000001111;
      patterns[721] = 50'b01_0000000000001011_0000000000000100_0000000000000111;
      patterns[722] = 50'b10_0000000000001011_0000000000000100_0000000000000000;
      patterns[723] = 50'b11_0000000000001011_0000000000000100_0000000000001111;
      patterns[724] = 50'b00_0000000000001011_0000000000000101_0000000000010000;
      patterns[725] = 50'b01_0000000000001011_0000000000000101_0000000000000110;
      patterns[726] = 50'b10_0000000000001011_0000000000000101_0000000000000001;
      patterns[727] = 50'b11_0000000000001011_0000000000000101_0000000000001111;
      patterns[728] = 50'b00_0000000000001011_0000000000000110_0000000000010001;
      patterns[729] = 50'b01_0000000000001011_0000000000000110_0000000000000101;
      patterns[730] = 50'b10_0000000000001011_0000000000000110_0000000000000010;
      patterns[731] = 50'b11_0000000000001011_0000000000000110_0000000000001111;
      patterns[732] = 50'b00_0000000000001011_0000000000000111_0000000000010010;
      patterns[733] = 50'b01_0000000000001011_0000000000000111_0000000000000100;
      patterns[734] = 50'b10_0000000000001011_0000000000000111_0000000000000011;
      patterns[735] = 50'b11_0000000000001011_0000000000000111_0000000000001111;
      patterns[736] = 50'b00_0000000000001011_0000000000001000_0000000000010011;
      patterns[737] = 50'b01_0000000000001011_0000000000001000_0000000000000011;
      patterns[738] = 50'b10_0000000000001011_0000000000001000_0000000000001000;
      patterns[739] = 50'b11_0000000000001011_0000000000001000_0000000000001011;
      patterns[740] = 50'b00_0000000000001011_0000000000001001_0000000000010100;
      patterns[741] = 50'b01_0000000000001011_0000000000001001_0000000000000010;
      patterns[742] = 50'b10_0000000000001011_0000000000001001_0000000000001001;
      patterns[743] = 50'b11_0000000000001011_0000000000001001_0000000000001011;
      patterns[744] = 50'b00_0000000000001011_0000000000001010_0000000000010101;
      patterns[745] = 50'b01_0000000000001011_0000000000001010_0000000000000001;
      patterns[746] = 50'b10_0000000000001011_0000000000001010_0000000000001010;
      patterns[747] = 50'b11_0000000000001011_0000000000001010_0000000000001011;
      patterns[748] = 50'b00_0000000000001011_0000000000001011_0000000000010110;
      patterns[749] = 50'b01_0000000000001011_0000000000001011_0000000000000000;
      patterns[750] = 50'b10_0000000000001011_0000000000001011_0000000000001011;
      patterns[751] = 50'b11_0000000000001011_0000000000001011_0000000000001011;
      patterns[752] = 50'b00_0000000000001011_0000000000001100_0000000000010111;
      patterns[753] = 50'b01_0000000000001011_0000000000001100_1111111111111111;
      patterns[754] = 50'b10_0000000000001011_0000000000001100_0000000000001000;
      patterns[755] = 50'b11_0000000000001011_0000000000001100_0000000000001111;
      patterns[756] = 50'b00_0000000000001011_0000000000001101_0000000000011000;
      patterns[757] = 50'b01_0000000000001011_0000000000001101_1111111111111110;
      patterns[758] = 50'b10_0000000000001011_0000000000001101_0000000000001001;
      patterns[759] = 50'b11_0000000000001011_0000000000001101_0000000000001111;
      patterns[760] = 50'b00_0000000000001011_0000000000001110_0000000000011001;
      patterns[761] = 50'b01_0000000000001011_0000000000001110_1111111111111101;
      patterns[762] = 50'b10_0000000000001011_0000000000001110_0000000000001010;
      patterns[763] = 50'b11_0000000000001011_0000000000001110_0000000000001111;
      patterns[764] = 50'b00_0000000000001011_0000000000001111_0000000000011010;
      patterns[765] = 50'b01_0000000000001011_0000000000001111_1111111111111100;
      patterns[766] = 50'b10_0000000000001011_0000000000001111_0000000000001011;
      patterns[767] = 50'b11_0000000000001011_0000000000001111_0000000000001111;
      patterns[768] = 50'b00_0000000000001100_0000000000000000_0000000000001100;
      patterns[769] = 50'b01_0000000000001100_0000000000000000_0000000000001100;
      patterns[770] = 50'b10_0000000000001100_0000000000000000_0000000000000000;
      patterns[771] = 50'b11_0000000000001100_0000000000000000_0000000000001100;
      patterns[772] = 50'b00_0000000000001100_0000000000000001_0000000000001101;
      patterns[773] = 50'b01_0000000000001100_0000000000000001_0000000000001011;
      patterns[774] = 50'b10_0000000000001100_0000000000000001_0000000000000000;
      patterns[775] = 50'b11_0000000000001100_0000000000000001_0000000000001101;
      patterns[776] = 50'b00_0000000000001100_0000000000000010_0000000000001110;
      patterns[777] = 50'b01_0000000000001100_0000000000000010_0000000000001010;
      patterns[778] = 50'b10_0000000000001100_0000000000000010_0000000000000000;
      patterns[779] = 50'b11_0000000000001100_0000000000000010_0000000000001110;
      patterns[780] = 50'b00_0000000000001100_0000000000000011_0000000000001111;
      patterns[781] = 50'b01_0000000000001100_0000000000000011_0000000000001001;
      patterns[782] = 50'b10_0000000000001100_0000000000000011_0000000000000000;
      patterns[783] = 50'b11_0000000000001100_0000000000000011_0000000000001111;
      patterns[784] = 50'b00_0000000000001100_0000000000000100_0000000000010000;
      patterns[785] = 50'b01_0000000000001100_0000000000000100_0000000000001000;
      patterns[786] = 50'b10_0000000000001100_0000000000000100_0000000000000100;
      patterns[787] = 50'b11_0000000000001100_0000000000000100_0000000000001100;
      patterns[788] = 50'b00_0000000000001100_0000000000000101_0000000000010001;
      patterns[789] = 50'b01_0000000000001100_0000000000000101_0000000000000111;
      patterns[790] = 50'b10_0000000000001100_0000000000000101_0000000000000100;
      patterns[791] = 50'b11_0000000000001100_0000000000000101_0000000000001101;
      patterns[792] = 50'b00_0000000000001100_0000000000000110_0000000000010010;
      patterns[793] = 50'b01_0000000000001100_0000000000000110_0000000000000110;
      patterns[794] = 50'b10_0000000000001100_0000000000000110_0000000000000100;
      patterns[795] = 50'b11_0000000000001100_0000000000000110_0000000000001110;
      patterns[796] = 50'b00_0000000000001100_0000000000000111_0000000000010011;
      patterns[797] = 50'b01_0000000000001100_0000000000000111_0000000000000101;
      patterns[798] = 50'b10_0000000000001100_0000000000000111_0000000000000100;
      patterns[799] = 50'b11_0000000000001100_0000000000000111_0000000000001111;
      patterns[800] = 50'b00_0000000000001100_0000000000001000_0000000000010100;
      patterns[801] = 50'b01_0000000000001100_0000000000001000_0000000000000100;
      patterns[802] = 50'b10_0000000000001100_0000000000001000_0000000000001000;
      patterns[803] = 50'b11_0000000000001100_0000000000001000_0000000000001100;
      patterns[804] = 50'b00_0000000000001100_0000000000001001_0000000000010101;
      patterns[805] = 50'b01_0000000000001100_0000000000001001_0000000000000011;
      patterns[806] = 50'b10_0000000000001100_0000000000001001_0000000000001000;
      patterns[807] = 50'b11_0000000000001100_0000000000001001_0000000000001101;
      patterns[808] = 50'b00_0000000000001100_0000000000001010_0000000000010110;
      patterns[809] = 50'b01_0000000000001100_0000000000001010_0000000000000010;
      patterns[810] = 50'b10_0000000000001100_0000000000001010_0000000000001000;
      patterns[811] = 50'b11_0000000000001100_0000000000001010_0000000000001110;
      patterns[812] = 50'b00_0000000000001100_0000000000001011_0000000000010111;
      patterns[813] = 50'b01_0000000000001100_0000000000001011_0000000000000001;
      patterns[814] = 50'b10_0000000000001100_0000000000001011_0000000000001000;
      patterns[815] = 50'b11_0000000000001100_0000000000001011_0000000000001111;
      patterns[816] = 50'b00_0000000000001100_0000000000001100_0000000000011000;
      patterns[817] = 50'b01_0000000000001100_0000000000001100_0000000000000000;
      patterns[818] = 50'b10_0000000000001100_0000000000001100_0000000000001100;
      patterns[819] = 50'b11_0000000000001100_0000000000001100_0000000000001100;
      patterns[820] = 50'b00_0000000000001100_0000000000001101_0000000000011001;
      patterns[821] = 50'b01_0000000000001100_0000000000001101_1111111111111111;
      patterns[822] = 50'b10_0000000000001100_0000000000001101_0000000000001100;
      patterns[823] = 50'b11_0000000000001100_0000000000001101_0000000000001101;
      patterns[824] = 50'b00_0000000000001100_0000000000001110_0000000000011010;
      patterns[825] = 50'b01_0000000000001100_0000000000001110_1111111111111110;
      patterns[826] = 50'b10_0000000000001100_0000000000001110_0000000000001100;
      patterns[827] = 50'b11_0000000000001100_0000000000001110_0000000000001110;
      patterns[828] = 50'b00_0000000000001100_0000000000001111_0000000000011011;
      patterns[829] = 50'b01_0000000000001100_0000000000001111_1111111111111101;
      patterns[830] = 50'b10_0000000000001100_0000000000001111_0000000000001100;
      patterns[831] = 50'b11_0000000000001100_0000000000001111_0000000000001111;
      patterns[832] = 50'b00_0000000000001101_0000000000000000_0000000000001101;
      patterns[833] = 50'b01_0000000000001101_0000000000000000_0000000000001101;
      patterns[834] = 50'b10_0000000000001101_0000000000000000_0000000000000000;
      patterns[835] = 50'b11_0000000000001101_0000000000000000_0000000000001101;
      patterns[836] = 50'b00_0000000000001101_0000000000000001_0000000000001110;
      patterns[837] = 50'b01_0000000000001101_0000000000000001_0000000000001100;
      patterns[838] = 50'b10_0000000000001101_0000000000000001_0000000000000001;
      patterns[839] = 50'b11_0000000000001101_0000000000000001_0000000000001101;
      patterns[840] = 50'b00_0000000000001101_0000000000000010_0000000000001111;
      patterns[841] = 50'b01_0000000000001101_0000000000000010_0000000000001011;
      patterns[842] = 50'b10_0000000000001101_0000000000000010_0000000000000000;
      patterns[843] = 50'b11_0000000000001101_0000000000000010_0000000000001111;
      patterns[844] = 50'b00_0000000000001101_0000000000000011_0000000000010000;
      patterns[845] = 50'b01_0000000000001101_0000000000000011_0000000000001010;
      patterns[846] = 50'b10_0000000000001101_0000000000000011_0000000000000001;
      patterns[847] = 50'b11_0000000000001101_0000000000000011_0000000000001111;
      patterns[848] = 50'b00_0000000000001101_0000000000000100_0000000000010001;
      patterns[849] = 50'b01_0000000000001101_0000000000000100_0000000000001001;
      patterns[850] = 50'b10_0000000000001101_0000000000000100_0000000000000100;
      patterns[851] = 50'b11_0000000000001101_0000000000000100_0000000000001101;
      patterns[852] = 50'b00_0000000000001101_0000000000000101_0000000000010010;
      patterns[853] = 50'b01_0000000000001101_0000000000000101_0000000000001000;
      patterns[854] = 50'b10_0000000000001101_0000000000000101_0000000000000101;
      patterns[855] = 50'b11_0000000000001101_0000000000000101_0000000000001101;
      patterns[856] = 50'b00_0000000000001101_0000000000000110_0000000000010011;
      patterns[857] = 50'b01_0000000000001101_0000000000000110_0000000000000111;
      patterns[858] = 50'b10_0000000000001101_0000000000000110_0000000000000100;
      patterns[859] = 50'b11_0000000000001101_0000000000000110_0000000000001111;
      patterns[860] = 50'b00_0000000000001101_0000000000000111_0000000000010100;
      patterns[861] = 50'b01_0000000000001101_0000000000000111_0000000000000110;
      patterns[862] = 50'b10_0000000000001101_0000000000000111_0000000000000101;
      patterns[863] = 50'b11_0000000000001101_0000000000000111_0000000000001111;
      patterns[864] = 50'b00_0000000000001101_0000000000001000_0000000000010101;
      patterns[865] = 50'b01_0000000000001101_0000000000001000_0000000000000101;
      patterns[866] = 50'b10_0000000000001101_0000000000001000_0000000000001000;
      patterns[867] = 50'b11_0000000000001101_0000000000001000_0000000000001101;
      patterns[868] = 50'b00_0000000000001101_0000000000001001_0000000000010110;
      patterns[869] = 50'b01_0000000000001101_0000000000001001_0000000000000100;
      patterns[870] = 50'b10_0000000000001101_0000000000001001_0000000000001001;
      patterns[871] = 50'b11_0000000000001101_0000000000001001_0000000000001101;
      patterns[872] = 50'b00_0000000000001101_0000000000001010_0000000000010111;
      patterns[873] = 50'b01_0000000000001101_0000000000001010_0000000000000011;
      patterns[874] = 50'b10_0000000000001101_0000000000001010_0000000000001000;
      patterns[875] = 50'b11_0000000000001101_0000000000001010_0000000000001111;
      patterns[876] = 50'b00_0000000000001101_0000000000001011_0000000000011000;
      patterns[877] = 50'b01_0000000000001101_0000000000001011_0000000000000010;
      patterns[878] = 50'b10_0000000000001101_0000000000001011_0000000000001001;
      patterns[879] = 50'b11_0000000000001101_0000000000001011_0000000000001111;
      patterns[880] = 50'b00_0000000000001101_0000000000001100_0000000000011001;
      patterns[881] = 50'b01_0000000000001101_0000000000001100_0000000000000001;
      patterns[882] = 50'b10_0000000000001101_0000000000001100_0000000000001100;
      patterns[883] = 50'b11_0000000000001101_0000000000001100_0000000000001101;
      patterns[884] = 50'b00_0000000000001101_0000000000001101_0000000000011010;
      patterns[885] = 50'b01_0000000000001101_0000000000001101_0000000000000000;
      patterns[886] = 50'b10_0000000000001101_0000000000001101_0000000000001101;
      patterns[887] = 50'b11_0000000000001101_0000000000001101_0000000000001101;
      patterns[888] = 50'b00_0000000000001101_0000000000001110_0000000000011011;
      patterns[889] = 50'b01_0000000000001101_0000000000001110_1111111111111111;
      patterns[890] = 50'b10_0000000000001101_0000000000001110_0000000000001100;
      patterns[891] = 50'b11_0000000000001101_0000000000001110_0000000000001111;
      patterns[892] = 50'b00_0000000000001101_0000000000001111_0000000000011100;
      patterns[893] = 50'b01_0000000000001101_0000000000001111_1111111111111110;
      patterns[894] = 50'b10_0000000000001101_0000000000001111_0000000000001101;
      patterns[895] = 50'b11_0000000000001101_0000000000001111_0000000000001111;
      patterns[896] = 50'b00_0000000000001110_0000000000000000_0000000000001110;
      patterns[897] = 50'b01_0000000000001110_0000000000000000_0000000000001110;
      patterns[898] = 50'b10_0000000000001110_0000000000000000_0000000000000000;
      patterns[899] = 50'b11_0000000000001110_0000000000000000_0000000000001110;
      patterns[900] = 50'b00_0000000000001110_0000000000000001_0000000000001111;
      patterns[901] = 50'b01_0000000000001110_0000000000000001_0000000000001101;
      patterns[902] = 50'b10_0000000000001110_0000000000000001_0000000000000000;
      patterns[903] = 50'b11_0000000000001110_0000000000000001_0000000000001111;
      patterns[904] = 50'b00_0000000000001110_0000000000000010_0000000000010000;
      patterns[905] = 50'b01_0000000000001110_0000000000000010_0000000000001100;
      patterns[906] = 50'b10_0000000000001110_0000000000000010_0000000000000010;
      patterns[907] = 50'b11_0000000000001110_0000000000000010_0000000000001110;
      patterns[908] = 50'b00_0000000000001110_0000000000000011_0000000000010001;
      patterns[909] = 50'b01_0000000000001110_0000000000000011_0000000000001011;
      patterns[910] = 50'b10_0000000000001110_0000000000000011_0000000000000010;
      patterns[911] = 50'b11_0000000000001110_0000000000000011_0000000000001111;
      patterns[912] = 50'b00_0000000000001110_0000000000000100_0000000000010010;
      patterns[913] = 50'b01_0000000000001110_0000000000000100_0000000000001010;
      patterns[914] = 50'b10_0000000000001110_0000000000000100_0000000000000100;
      patterns[915] = 50'b11_0000000000001110_0000000000000100_0000000000001110;
      patterns[916] = 50'b00_0000000000001110_0000000000000101_0000000000010011;
      patterns[917] = 50'b01_0000000000001110_0000000000000101_0000000000001001;
      patterns[918] = 50'b10_0000000000001110_0000000000000101_0000000000000100;
      patterns[919] = 50'b11_0000000000001110_0000000000000101_0000000000001111;
      patterns[920] = 50'b00_0000000000001110_0000000000000110_0000000000010100;
      patterns[921] = 50'b01_0000000000001110_0000000000000110_0000000000001000;
      patterns[922] = 50'b10_0000000000001110_0000000000000110_0000000000000110;
      patterns[923] = 50'b11_0000000000001110_0000000000000110_0000000000001110;
      patterns[924] = 50'b00_0000000000001110_0000000000000111_0000000000010101;
      patterns[925] = 50'b01_0000000000001110_0000000000000111_0000000000000111;
      patterns[926] = 50'b10_0000000000001110_0000000000000111_0000000000000110;
      patterns[927] = 50'b11_0000000000001110_0000000000000111_0000000000001111;
      patterns[928] = 50'b00_0000000000001110_0000000000001000_0000000000010110;
      patterns[929] = 50'b01_0000000000001110_0000000000001000_0000000000000110;
      patterns[930] = 50'b10_0000000000001110_0000000000001000_0000000000001000;
      patterns[931] = 50'b11_0000000000001110_0000000000001000_0000000000001110;
      patterns[932] = 50'b00_0000000000001110_0000000000001001_0000000000010111;
      patterns[933] = 50'b01_0000000000001110_0000000000001001_0000000000000101;
      patterns[934] = 50'b10_0000000000001110_0000000000001001_0000000000001000;
      patterns[935] = 50'b11_0000000000001110_0000000000001001_0000000000001111;
      patterns[936] = 50'b00_0000000000001110_0000000000001010_0000000000011000;
      patterns[937] = 50'b01_0000000000001110_0000000000001010_0000000000000100;
      patterns[938] = 50'b10_0000000000001110_0000000000001010_0000000000001010;
      patterns[939] = 50'b11_0000000000001110_0000000000001010_0000000000001110;
      patterns[940] = 50'b00_0000000000001110_0000000000001011_0000000000011001;
      patterns[941] = 50'b01_0000000000001110_0000000000001011_0000000000000011;
      patterns[942] = 50'b10_0000000000001110_0000000000001011_0000000000001010;
      patterns[943] = 50'b11_0000000000001110_0000000000001011_0000000000001111;
      patterns[944] = 50'b00_0000000000001110_0000000000001100_0000000000011010;
      patterns[945] = 50'b01_0000000000001110_0000000000001100_0000000000000010;
      patterns[946] = 50'b10_0000000000001110_0000000000001100_0000000000001100;
      patterns[947] = 50'b11_0000000000001110_0000000000001100_0000000000001110;
      patterns[948] = 50'b00_0000000000001110_0000000000001101_0000000000011011;
      patterns[949] = 50'b01_0000000000001110_0000000000001101_0000000000000001;
      patterns[950] = 50'b10_0000000000001110_0000000000001101_0000000000001100;
      patterns[951] = 50'b11_0000000000001110_0000000000001101_0000000000001111;
      patterns[952] = 50'b00_0000000000001110_0000000000001110_0000000000011100;
      patterns[953] = 50'b01_0000000000001110_0000000000001110_0000000000000000;
      patterns[954] = 50'b10_0000000000001110_0000000000001110_0000000000001110;
      patterns[955] = 50'b11_0000000000001110_0000000000001110_0000000000001110;
      patterns[956] = 50'b00_0000000000001110_0000000000001111_0000000000011101;
      patterns[957] = 50'b01_0000000000001110_0000000000001111_1111111111111111;
      patterns[958] = 50'b10_0000000000001110_0000000000001111_0000000000001110;
      patterns[959] = 50'b11_0000000000001110_0000000000001111_0000000000001111;
      patterns[960] = 50'b00_0000000000001111_0000000000000000_0000000000001111;
      patterns[961] = 50'b01_0000000000001111_0000000000000000_0000000000001111;
      patterns[962] = 50'b10_0000000000001111_0000000000000000_0000000000000000;
      patterns[963] = 50'b11_0000000000001111_0000000000000000_0000000000001111;
      patterns[964] = 50'b00_0000000000001111_0000000000000001_0000000000010000;
      patterns[965] = 50'b01_0000000000001111_0000000000000001_0000000000001110;
      patterns[966] = 50'b10_0000000000001111_0000000000000001_0000000000000001;
      patterns[967] = 50'b11_0000000000001111_0000000000000001_0000000000001111;
      patterns[968] = 50'b00_0000000000001111_0000000000000010_0000000000010001;
      patterns[969] = 50'b01_0000000000001111_0000000000000010_0000000000001101;
      patterns[970] = 50'b10_0000000000001111_0000000000000010_0000000000000010;
      patterns[971] = 50'b11_0000000000001111_0000000000000010_0000000000001111;
      patterns[972] = 50'b00_0000000000001111_0000000000000011_0000000000010010;
      patterns[973] = 50'b01_0000000000001111_0000000000000011_0000000000001100;
      patterns[974] = 50'b10_0000000000001111_0000000000000011_0000000000000011;
      patterns[975] = 50'b11_0000000000001111_0000000000000011_0000000000001111;
      patterns[976] = 50'b00_0000000000001111_0000000000000100_0000000000010011;
      patterns[977] = 50'b01_0000000000001111_0000000000000100_0000000000001011;
      patterns[978] = 50'b10_0000000000001111_0000000000000100_0000000000000100;
      patterns[979] = 50'b11_0000000000001111_0000000000000100_0000000000001111;
      patterns[980] = 50'b00_0000000000001111_0000000000000101_0000000000010100;
      patterns[981] = 50'b01_0000000000001111_0000000000000101_0000000000001010;
      patterns[982] = 50'b10_0000000000001111_0000000000000101_0000000000000101;
      patterns[983] = 50'b11_0000000000001111_0000000000000101_0000000000001111;
      patterns[984] = 50'b00_0000000000001111_0000000000000110_0000000000010101;
      patterns[985] = 50'b01_0000000000001111_0000000000000110_0000000000001001;
      patterns[986] = 50'b10_0000000000001111_0000000000000110_0000000000000110;
      patterns[987] = 50'b11_0000000000001111_0000000000000110_0000000000001111;
      patterns[988] = 50'b00_0000000000001111_0000000000000111_0000000000010110;
      patterns[989] = 50'b01_0000000000001111_0000000000000111_0000000000001000;
      patterns[990] = 50'b10_0000000000001111_0000000000000111_0000000000000111;
      patterns[991] = 50'b11_0000000000001111_0000000000000111_0000000000001111;
      patterns[992] = 50'b00_0000000000001111_0000000000001000_0000000000010111;
      patterns[993] = 50'b01_0000000000001111_0000000000001000_0000000000000111;
      patterns[994] = 50'b10_0000000000001111_0000000000001000_0000000000001000;
      patterns[995] = 50'b11_0000000000001111_0000000000001000_0000000000001111;
      patterns[996] = 50'b00_0000000000001111_0000000000001001_0000000000011000;
      patterns[997] = 50'b01_0000000000001111_0000000000001001_0000000000000110;
      patterns[998] = 50'b10_0000000000001111_0000000000001001_0000000000001001;
      patterns[999] = 50'b11_0000000000001111_0000000000001001_0000000000001111;
      patterns[1000] = 50'b00_0000000000001111_0000000000001010_0000000000011001;
      patterns[1001] = 50'b01_0000000000001111_0000000000001010_0000000000000101;
      patterns[1002] = 50'b10_0000000000001111_0000000000001010_0000000000001010;
      patterns[1003] = 50'b11_0000000000001111_0000000000001010_0000000000001111;
      patterns[1004] = 50'b00_0000000000001111_0000000000001011_0000000000011010;
      patterns[1005] = 50'b01_0000000000001111_0000000000001011_0000000000000100;
      patterns[1006] = 50'b10_0000000000001111_0000000000001011_0000000000001011;
      patterns[1007] = 50'b11_0000000000001111_0000000000001011_0000000000001111;
      patterns[1008] = 50'b00_0000000000001111_0000000000001100_0000000000011011;
      patterns[1009] = 50'b01_0000000000001111_0000000000001100_0000000000000011;
      patterns[1010] = 50'b10_0000000000001111_0000000000001100_0000000000001100;
      patterns[1011] = 50'b11_0000000000001111_0000000000001100_0000000000001111;
      patterns[1012] = 50'b00_0000000000001111_0000000000001101_0000000000011100;
      patterns[1013] = 50'b01_0000000000001111_0000000000001101_0000000000000010;
      patterns[1014] = 50'b10_0000000000001111_0000000000001101_0000000000001101;
      patterns[1015] = 50'b11_0000000000001111_0000000000001101_0000000000001111;
      patterns[1016] = 50'b00_0000000000001111_0000000000001110_0000000000011101;
      patterns[1017] = 50'b01_0000000000001111_0000000000001110_0000000000000001;
      patterns[1018] = 50'b10_0000000000001111_0000000000001110_0000000000001110;
      patterns[1019] = 50'b11_0000000000001111_0000000000001110_0000000000001111;
      patterns[1020] = 50'b00_0000000000001111_0000000000001111_0000000000011110;
      patterns[1021] = 50'b01_0000000000001111_0000000000001111_0000000000000000;
      patterns[1022] = 50'b10_0000000000001111_0000000000001111_0000000000001111;
      patterns[1023] = 50'b11_0000000000001111_0000000000001111_0000000000001111;
      patterns[1024] = 50'b00_1101111011101000_0111000010100000_0100111110001000;
      patterns[1025] = 50'b01_1101111011101000_0111000010100000_0110111001001000;
      patterns[1026] = 50'b10_1101111011101000_0111000010100000_0101000010100000;
      patterns[1027] = 50'b11_1101111011101000_0111000010100000_1111111011101000;
      patterns[1028] = 50'b00_1001011111010011_0010010001101000_1011110000111011;
      patterns[1029] = 50'b01_1001011111010011_0010010001101000_0111001101101011;
      patterns[1030] = 50'b10_1001011111010011_0010010001101000_0000010001000000;
      patterns[1031] = 50'b11_1001011111010011_0010010001101000_1011011111111011;
      patterns[1032] = 50'b00_1000000101100101_0111111010110010_0000000000010111;
      patterns[1033] = 50'b01_1000000101100101_0111111010110010_0000001010110011;
      patterns[1034] = 50'b10_1000000101100101_0111111010110010_0000000000100000;
      patterns[1035] = 50'b11_1000000101100101_0111111010110010_1111111111110111;
      patterns[1036] = 50'b00_1001100100110011_0011100000111010_1101000101101101;
      patterns[1037] = 50'b01_1001100100110011_0011100000111010_0110000011111001;
      patterns[1038] = 50'b10_1001100100110011_0011100000111010_0001100000110010;
      patterns[1039] = 50'b11_1001100100110011_0011100000111010_1011100100111011;
      patterns[1040] = 50'b00_1101001000100101_0011100001001111_0000101001110100;
      patterns[1041] = 50'b01_1101001000100101_0011100001001111_1001100111010110;
      patterns[1042] = 50'b10_1101001000100101_0011100001001111_0001000000000101;
      patterns[1043] = 50'b11_1101001000100101_0011100001001111_1111101001101111;
      patterns[1044] = 50'b00_0001000011110100_1111000100000000_0000000111110100;
      patterns[1045] = 50'b01_0001000011110100_1111000100000000_0001111111110100;
      patterns[1046] = 50'b10_0001000011110100_1111000100000000_0001000000000000;
      patterns[1047] = 50'b11_0001000011110100_1111000100000000_1111000111110100;
      patterns[1048] = 50'b00_0110110001111010_0011011001111100_1010001011110110;
      patterns[1049] = 50'b01_0110110001111010_0011011001111100_0011010111111110;
      patterns[1050] = 50'b10_0110110001111010_0011011001111100_0010010001111000;
      patterns[1051] = 50'b11_0110110001111010_0011011001111100_0111111001111110;
      patterns[1052] = 50'b00_1110000110000100_1001101011001000_0111110001001100;
      patterns[1053] = 50'b01_1110000110000100_1001101011001000_0100011010111100;
      patterns[1054] = 50'b10_1110000110000100_1001101011001000_1000000010000000;
      patterns[1055] = 50'b11_1110000110000100_1001101011001000_1111101111001100;
      patterns[1056] = 50'b00_0111001100101011_1111100001001000_0110101101110011;
      patterns[1057] = 50'b01_0111001100101011_1111100001001000_0111101011100011;
      patterns[1058] = 50'b10_0111001100101011_1111100001001000_0111000000001000;
      patterns[1059] = 50'b11_0111001100101011_1111100001001000_1111101101101011;
      patterns[1060] = 50'b00_1110011000110011_1100011111110110_1010111000101001;
      patterns[1061] = 50'b01_1110011000110011_1100011111110110_0001111000111101;
      patterns[1062] = 50'b10_1110011000110011_1100011111110110_1100011000110010;
      patterns[1063] = 50'b11_1110011000110011_1100011111110110_1110011111110111;
      patterns[1064] = 50'b00_1001110110101001_1111101000011110_1001011111000111;
      patterns[1065] = 50'b01_1001110110101001_1111101000011110_1010001110001011;
      patterns[1066] = 50'b10_1001110110101001_1111101000011110_1001100000001000;
      patterns[1067] = 50'b11_1001110110101001_1111101000011110_1111111110111111;
      patterns[1068] = 50'b00_0110000101011010_0101010111111011_1011011101010101;
      patterns[1069] = 50'b01_0110000101011010_0101010111111011_0000101101011111;
      patterns[1070] = 50'b10_0110000101011010_0101010111111011_0100000101011010;
      patterns[1071] = 50'b11_0110000101011010_0101010111111011_0111010111111011;
      patterns[1072] = 50'b00_0010000111101010_0110010001000101_1000011000101111;
      patterns[1073] = 50'b01_0010000111101010_0110010001000101_1011110110100101;
      patterns[1074] = 50'b10_0010000111101010_0110010001000101_0010000001000000;
      patterns[1075] = 50'b11_0010000111101010_0110010001000101_0110010111101111;
      patterns[1076] = 50'b00_1101001010010000_1100111001000001_1010000011010001;
      patterns[1077] = 50'b01_1101001010010000_1100111001000001_0000010001001111;
      patterns[1078] = 50'b10_1101001010010000_1100111001000001_1100001000000000;
      patterns[1079] = 50'b11_1101001010010000_1100111001000001_1101111011010001;
      patterns[1080] = 50'b00_1011010000010000_0000110101110111_1100000110000111;
      patterns[1081] = 50'b01_1011010000010000_0000110101110111_1010011010011001;
      patterns[1082] = 50'b10_1011010000010000_0000110101110111_0000010000010000;
      patterns[1083] = 50'b11_1011010000010000_0000110101110111_1011110101110111;
      patterns[1084] = 50'b00_1000011111001000_1010001010111101_0010101010000101;
      patterns[1085] = 50'b01_1000011111001000_1010001010111101_1110010100001011;
      patterns[1086] = 50'b10_1000011111001000_1010001010111101_1000001010001000;
      patterns[1087] = 50'b11_1000011111001000_1010001010111101_1010011111111101;
      patterns[1088] = 50'b00_0000001001101011_1001110101111011_1001111111100110;
      patterns[1089] = 50'b01_0000001001101011_1001110101111011_0110010011110000;
      patterns[1090] = 50'b10_0000001001101011_1001110101111011_0000000001101011;
      patterns[1091] = 50'b11_0000001001101011_1001110101111011_1001111101111011;
      patterns[1092] = 50'b00_1111110101111010_1000100011010001_1000011001001011;
      patterns[1093] = 50'b01_1111110101111010_1000100011010001_0111010010101001;
      patterns[1094] = 50'b10_1111110101111010_1000100011010001_1000100001010000;
      patterns[1095] = 50'b11_1111110101111010_1000100011010001_1111110111111011;
      patterns[1096] = 50'b00_1010100101110111_0101001100100000_1111110010010111;
      patterns[1097] = 50'b01_1010100101110111_0101001100100000_0101011001010111;
      patterns[1098] = 50'b10_1010100101110111_0101001100100000_0000000100100000;
      patterns[1099] = 50'b11_1010100101110111_0101001100100000_1111101101110111;
      patterns[1100] = 50'b00_1100101100101010_0010000001100000_1110101110001010;
      patterns[1101] = 50'b01_1100101100101010_0010000001100000_1010101011001010;
      patterns[1102] = 50'b10_1100101100101010_0010000001100000_0000000000100000;
      patterns[1103] = 50'b11_1100101100101010_0010000001100000_1110101101101010;
      patterns[1104] = 50'b00_1001100011101101_0101000000100001_1110100100001110;
      patterns[1105] = 50'b01_1001100011101101_0101000000100001_0100100011001100;
      patterns[1106] = 50'b10_1001100011101101_0101000000100001_0001000000100001;
      patterns[1107] = 50'b11_1001100011101101_0101000000100001_1101100011101101;
      patterns[1108] = 50'b00_0110101011100000_0010100001001100_1001001100101100;
      patterns[1109] = 50'b01_0110101011100000_0010100001001100_0100001010010100;
      patterns[1110] = 50'b10_0110101011100000_0010100001001100_0010100001000000;
      patterns[1111] = 50'b11_0110101011100000_0010100001001100_0110101011101100;
      patterns[1112] = 50'b00_0100100000001100_0101010010101101_1001110010111001;
      patterns[1113] = 50'b01_0100100000001100_0101010010101101_1111001101011111;
      patterns[1114] = 50'b10_0100100000001100_0101010010101101_0100000000001100;
      patterns[1115] = 50'b11_0100100000001100_0101010010101101_0101110010101101;
      patterns[1116] = 50'b00_1010001101111110_1011110010111000_0110000000110110;
      patterns[1117] = 50'b01_1010001101111110_1011110010111000_1110011011000110;
      patterns[1118] = 50'b10_1010001101111110_1011110010111000_1010000000111000;
      patterns[1119] = 50'b11_1010001101111110_1011110010111000_1011111111111110;
      patterns[1120] = 50'b00_1110010010010111_1000001110110000_0110100001000111;
      patterns[1121] = 50'b01_1110010010010111_1000001110110000_0110000011100111;
      patterns[1122] = 50'b10_1110010010010111_1000001110110000_1000000010010000;
      patterns[1123] = 50'b11_1110010010010111_1000001110110000_1110011110110111;
      patterns[1124] = 50'b00_1011111100000001_0111111011000011_0011110111000100;
      patterns[1125] = 50'b01_1011111100000001_0111111011000011_0100000000111110;
      patterns[1126] = 50'b10_1011111100000001_0111111011000011_0011111000000001;
      patterns[1127] = 50'b11_1011111100000001_0111111011000011_1111111111000011;
      patterns[1128] = 50'b00_1101110101001000_0010000000100000_1111110101101000;
      patterns[1129] = 50'b01_1101110101001000_0010000000100000_1011110100101000;
      patterns[1130] = 50'b10_1101110101001000_0010000000100000_0000000000000000;
      patterns[1131] = 50'b11_1101110101001000_0010000000100000_1111110101101000;
      patterns[1132] = 50'b00_1111111100000100_0001000010100101_0000111110101001;
      patterns[1133] = 50'b01_1111111100000100_0001000010100101_1110111001011111;
      patterns[1134] = 50'b10_1111111100000100_0001000010100101_0001000000000100;
      patterns[1135] = 50'b11_1111111100000100_0001000010100101_1111111110100101;
      patterns[1136] = 50'b00_1100010110110110_0011001011001110_1111100010000100;
      patterns[1137] = 50'b01_1100010110110110_0011001011001110_1001001011101000;
      patterns[1138] = 50'b10_1100010110110110_0011001011001110_0000000010000110;
      patterns[1139] = 50'b11_1100010110110110_0011001011001110_1111011111111110;
      patterns[1140] = 50'b00_1111001100101001_0000010001010011_1111011101111100;
      patterns[1141] = 50'b01_1111001100101001_0000010001010011_1110111011010110;
      patterns[1142] = 50'b10_1111001100101001_0000010001010011_0000000000000001;
      patterns[1143] = 50'b11_1111001100101001_0000010001010011_1111011101111011;
      patterns[1144] = 50'b00_1001011011010011_1010111110011010_0100011001101101;
      patterns[1145] = 50'b01_1001011011010011_1010111110011010_1110011100111001;
      patterns[1146] = 50'b10_1001011011010011_1010111110011010_1000011010010010;
      patterns[1147] = 50'b11_1001011011010011_1010111110011010_1011111111011011;
      patterns[1148] = 50'b00_0110111000111101_0011011000010110_1010010001010011;
      patterns[1149] = 50'b01_0110111000111101_0011011000010110_0011100000100111;
      patterns[1150] = 50'b10_0110111000111101_0011011000010110_0010011000010100;
      patterns[1151] = 50'b11_0110111000111101_0011011000010110_0111111000111111;
      patterns[1152] = 50'b00_1011110010011011_1111111111111001_1011110010010100;
      patterns[1153] = 50'b01_1011110010011011_1111111111111001_1011110010100010;
      patterns[1154] = 50'b10_1011110010011011_1111111111111001_1011110010011001;
      patterns[1155] = 50'b11_1011110010011011_1111111111111001_1111111111111011;
      patterns[1156] = 50'b00_1101100000101111_1000111111000010_0110011111110001;
      patterns[1157] = 50'b01_1101100000101111_1000111111000010_0100100001101101;
      patterns[1158] = 50'b10_1101100000101111_1000111111000010_1000100000000010;
      patterns[1159] = 50'b11_1101100000101111_1000111111000010_1101111111101111;
      patterns[1160] = 50'b00_0011011010001100_1101000000110100_0000011011000000;
      patterns[1161] = 50'b01_0011011010001100_1101000000110100_0110011001011000;
      patterns[1162] = 50'b10_0011011010001100_1101000000110100_0001000000000100;
      patterns[1163] = 50'b11_0011011010001100_1101000000110100_1111011010111100;
      patterns[1164] = 50'b00_1000010000111000_0101110001110110_1110000010101110;
      patterns[1165] = 50'b01_1000010000111000_0101110001110110_0010011111000010;
      patterns[1166] = 50'b10_1000010000111000_0101110001110110_0000010000110000;
      patterns[1167] = 50'b11_1000010000111000_0101110001110110_1101110001111110;
      patterns[1168] = 50'b00_0100111000000100_1001101111010110_1110100111011010;
      patterns[1169] = 50'b01_0100111000000100_1001101111010110_1011001000101110;
      patterns[1170] = 50'b10_0100111000000100_1001101111010110_0000101000000100;
      patterns[1171] = 50'b11_0100111000000100_1001101111010110_1101111111010110;
      patterns[1172] = 50'b00_1000001111001110_1010100000001010_0010101111011000;
      patterns[1173] = 50'b01_1000001111001110_1010100000001010_1101101111000100;
      patterns[1174] = 50'b10_1000001111001110_1010100000001010_1000000000001010;
      patterns[1175] = 50'b11_1000001111001110_1010100000001010_1010101111001110;
      patterns[1176] = 50'b00_0000101010011100_1011110100010101_1100011110110001;
      patterns[1177] = 50'b01_0000101010011100_1011110100010101_0100110110000111;
      patterns[1178] = 50'b10_0000101010011100_1011110100010101_0000100000010100;
      patterns[1179] = 50'b11_0000101010011100_1011110100010101_1011111110011101;
      patterns[1180] = 50'b00_0010100000110110_1010000010011010_1100100011010000;
      patterns[1181] = 50'b01_0010100000110110_1010000010011010_1000011110011100;
      patterns[1182] = 50'b10_0010100000110110_1010000010011010_0010000000010010;
      patterns[1183] = 50'b11_0010100000110110_1010000010011010_1010100010111110;
      patterns[1184] = 50'b00_1001101000011011_1011001001001000_0100110001100011;
      patterns[1185] = 50'b01_1001101000011011_1011001001001000_1110011111010011;
      patterns[1186] = 50'b10_1001101000011011_1011001001001000_1001001000001000;
      patterns[1187] = 50'b11_1001101000011011_1011001001001000_1011101001011011;
      patterns[1188] = 50'b00_0000010111010101_1001001111011010_1001100110101111;
      patterns[1189] = 50'b01_0000010111010101_1001001111011010_0111000111111011;
      patterns[1190] = 50'b10_0000010111010101_1001001111011010_0000000111010000;
      patterns[1191] = 50'b11_0000010111010101_1001001111011010_1001011111011111;
      patterns[1192] = 50'b00_0101011010100001_1110001110110100_0011101001010101;
      patterns[1193] = 50'b01_0101011010100001_1110001110110100_0111001011101101;
      patterns[1194] = 50'b10_0101011010100001_1110001110110100_0100001010100000;
      patterns[1195] = 50'b11_0101011010100001_1110001110110100_1111011110110101;
      patterns[1196] = 50'b00_1101010110011110_1110110100010111_1100001010110101;
      patterns[1197] = 50'b01_1101010110011110_1110110100010111_1110100010000111;
      patterns[1198] = 50'b10_1101010110011110_1110110100010111_1100010100010110;
      patterns[1199] = 50'b11_1101010110011110_1110110100010111_1111110110011111;
      patterns[1200] = 50'b00_1111001100001110_0111001100101001_0110011000110111;
      patterns[1201] = 50'b01_1111001100001110_0111001100101001_0111111111100101;
      patterns[1202] = 50'b10_1111001100001110_0111001100101001_0111001100001000;
      patterns[1203] = 50'b11_1111001100001110_0111001100101001_1111001100101111;
      patterns[1204] = 50'b00_0000001000100110_1000110000001111_1000111000110101;
      patterns[1205] = 50'b01_0000001000100110_1000110000001111_0111011000010111;
      patterns[1206] = 50'b10_0000001000100110_1000110000001111_0000000000000110;
      patterns[1207] = 50'b11_0000001000100110_1000110000001111_1000111000101111;
      patterns[1208] = 50'b00_1001101011101010_1000011001010110_0010000101000000;
      patterns[1209] = 50'b01_1001101011101010_1000011001010110_0001010010010100;
      patterns[1210] = 50'b10_1001101011101010_1000011001010110_1000001001000010;
      patterns[1211] = 50'b11_1001101011101010_1000011001010110_1001111011111110;
      patterns[1212] = 50'b00_0000011101001101_1110100000010100_1110111101100001;
      patterns[1213] = 50'b01_0000011101001101_1110100000010100_0001111100111001;
      patterns[1214] = 50'b10_0000011101001101_1110100000010100_0000000000000100;
      patterns[1215] = 50'b11_0000011101001101_1110100000010100_1110111101011101;
      patterns[1216] = 50'b00_1000000000110000_0000101110111111_1000101111101111;
      patterns[1217] = 50'b01_1000000000110000_0000101110111111_0111010001110001;
      patterns[1218] = 50'b10_1000000000110000_0000101110111111_0000000000110000;
      patterns[1219] = 50'b11_1000000000110000_0000101110111111_1000101110111111;
      patterns[1220] = 50'b00_0000110010001010_1011011000010111_1100001010100001;
      patterns[1221] = 50'b01_0000110010001010_1011011000010111_0101011001110011;
      patterns[1222] = 50'b10_0000110010001010_1011011000010111_0000010000000010;
      patterns[1223] = 50'b11_0000110010001010_1011011000010111_1011111010011111;
      patterns[1224] = 50'b00_0110011011001100_0011000110111011_1001100010000111;
      patterns[1225] = 50'b01_0110011011001100_0011000110111011_0011010100010001;
      patterns[1226] = 50'b10_0110011011001100_0011000110111011_0010000010001000;
      patterns[1227] = 50'b11_0110011011001100_0011000110111011_0111011111111111;
      patterns[1228] = 50'b00_0100101100110001_0011001110001101_0111111010111110;
      patterns[1229] = 50'b01_0100101100110001_0011001110001101_0001011110100100;
      patterns[1230] = 50'b10_0100101100110001_0011001110001101_0000001100000001;
      patterns[1231] = 50'b11_0100101100110001_0011001110001101_0111101110111101;
      patterns[1232] = 50'b00_0011101010111011_1010010111101000_1110000010100011;
      patterns[1233] = 50'b01_0011101010111011_1010010111101000_1001010011010011;
      patterns[1234] = 50'b10_0011101010111011_1010010111101000_0010000010101000;
      patterns[1235] = 50'b11_0011101010111011_1010010111101000_1011111111111011;
      patterns[1236] = 50'b00_1110001101011010_1100101101010101_1010111010101111;
      patterns[1237] = 50'b01_1110001101011010_1100101101010101_0001100000000101;
      patterns[1238] = 50'b10_1110001101011010_1100101101010101_1100001101010000;
      patterns[1239] = 50'b11_1110001101011010_1100101101010101_1110101101011111;
      patterns[1240] = 50'b00_1010001100000110_0011101100000000_1101111000000110;
      patterns[1241] = 50'b01_1010001100000110_0011101100000000_0110100000000110;
      patterns[1242] = 50'b10_1010001100000110_0011101100000000_0010001100000000;
      patterns[1243] = 50'b11_1010001100000110_0011101100000000_1011101100000110;
      patterns[1244] = 50'b00_1011101100111001_1000010100001010_0100000001000011;
      patterns[1245] = 50'b01_1011101100111001_1000010100001010_0011011000101111;
      patterns[1246] = 50'b10_1011101100111001_1000010100001010_1000000100001000;
      patterns[1247] = 50'b11_1011101100111001_1000010100001010_1011111100111011;
      patterns[1248] = 50'b00_1101000100011100_1100000111110100_1001001100010000;
      patterns[1249] = 50'b01_1101000100011100_1100000111110100_0000111100101000;
      patterns[1250] = 50'b10_1101000100011100_1100000111110100_1100000100010100;
      patterns[1251] = 50'b11_1101000100011100_1100000111110100_1101000111111100;
      patterns[1252] = 50'b00_1110010111111111_1001001001101101_0111100001101100;
      patterns[1253] = 50'b01_1110010111111111_1001001001101101_0101001110010010;
      patterns[1254] = 50'b10_1110010111111111_1001001001101101_1000000001101101;
      patterns[1255] = 50'b11_1110010111111111_1001001001101101_1111011111111111;
      patterns[1256] = 50'b00_1000000100111000_1011101010110111_0011101111101111;
      patterns[1257] = 50'b01_1000000100111000_1011101010110111_1100011010000001;
      patterns[1258] = 50'b10_1000000100111000_1011101010110111_1000000000110000;
      patterns[1259] = 50'b11_1000000100111000_1011101010110111_1011101110111111;
      patterns[1260] = 50'b00_1101100010100101_0101100111001011_0011001001110000;
      patterns[1261] = 50'b01_1101100010100101_0101100111001011_0111111011011010;
      patterns[1262] = 50'b10_1101100010100101_0101100111001011_0101100010000001;
      patterns[1263] = 50'b11_1101100010100101_0101100111001011_1101100111101111;
      patterns[1264] = 50'b00_0011110111011001_0000000000110010_0011111000001011;
      patterns[1265] = 50'b01_0011110111011001_0000000000110010_0011110110100111;
      patterns[1266] = 50'b10_0011110111011001_0000000000110010_0000000000010000;
      patterns[1267] = 50'b11_0011110111011001_0000000000110010_0011110111111011;
      patterns[1268] = 50'b00_0110010000111101_1000111110001110_1111001111001011;
      patterns[1269] = 50'b01_0110010000111101_1000111110001110_1101010010101111;
      patterns[1270] = 50'b10_0110010000111101_1000111110001110_0000010000001100;
      patterns[1271] = 50'b11_0110010000111101_1000111110001110_1110111110111111;
      patterns[1272] = 50'b00_0111110101111000_1011101000101110_0011011110100110;
      patterns[1273] = 50'b01_0111110101111000_1011101000101110_1100001101001010;
      patterns[1274] = 50'b10_0111110101111000_1011101000101110_0011100000101000;
      patterns[1275] = 50'b11_0111110101111000_1011101000101110_1111111101111110;
      patterns[1276] = 50'b00_0000011010010111_0100110001100101_0101001011111100;
      patterns[1277] = 50'b01_0000011010010111_0100110001100101_1011101000110010;
      patterns[1278] = 50'b10_0000011010010111_0100110001100101_0000010000000101;
      patterns[1279] = 50'b11_0000011010010111_0100110001100101_0100111011110111;
      patterns[1280] = 50'b00_0001111100001000_1010111100111100_1100111001000100;
      patterns[1281] = 50'b01_0001111100001000_1010111100111100_0110111111001100;
      patterns[1282] = 50'b10_0001111100001000_1010111100111100_0000111100001000;
      patterns[1283] = 50'b11_0001111100001000_1010111100111100_1011111100111100;
      patterns[1284] = 50'b00_1010001101011111_1001000010100110_0011010000000101;
      patterns[1285] = 50'b01_1010001101011111_1001000010100110_0001001010111001;
      patterns[1286] = 50'b10_1010001101011111_1001000010100110_1000000000000110;
      patterns[1287] = 50'b11_1010001101011111_1001000010100110_1011001111111111;
      patterns[1288] = 50'b00_0001111011101011_1000011111110001_1010011011011100;
      patterns[1289] = 50'b01_0001111011101011_1000011111110001_1001011011111010;
      patterns[1290] = 50'b10_0001111011101011_1000011111110001_0000011011100001;
      patterns[1291] = 50'b11_0001111011101011_1000011111110001_1001111111111011;
      patterns[1292] = 50'b00_0010000100001000_0101000011011001_0111000111100001;
      patterns[1293] = 50'b01_0010000100001000_0101000011011001_1101000000101111;
      patterns[1294] = 50'b10_0010000100001000_0101000011011001_0000000000001000;
      patterns[1295] = 50'b11_0010000100001000_0101000011011001_0111000111011001;
      patterns[1296] = 50'b00_0001101101011011_1011001111101001_1100111101000100;
      patterns[1297] = 50'b01_0001101101011011_1011001111101001_0110011101110010;
      patterns[1298] = 50'b10_0001101101011011_1011001111101001_0001001101001001;
      patterns[1299] = 50'b11_0001101101011011_1011001111101001_1011101111111011;
      patterns[1300] = 50'b00_1011011000100111_1111101010010101_1011000010111100;
      patterns[1301] = 50'b01_1011011000100111_1111101010010101_1011101110010010;
      patterns[1302] = 50'b10_1011011000100111_1111101010010101_1011001000000101;
      patterns[1303] = 50'b11_1011011000100111_1111101010010101_1111111010110111;
      patterns[1304] = 50'b00_0110010010000011_0110100001111001_1100110011111100;
      patterns[1305] = 50'b01_0110010010000011_0110100001111001_1111110000001010;
      patterns[1306] = 50'b10_0110010010000011_0110100001111001_0110000000000001;
      patterns[1307] = 50'b11_0110010010000011_0110100001111001_0110110011111011;
      patterns[1308] = 50'b00_1110110100001000_0101110000011000_0100100100100000;
      patterns[1309] = 50'b01_1110110100001000_0101110000011000_1001000011110000;
      patterns[1310] = 50'b10_1110110100001000_0101110000011000_0100110000001000;
      patterns[1311] = 50'b11_1110110100001000_0101110000011000_1111110100011000;
      patterns[1312] = 50'b00_1110000110111111_1001111111111011_1000000110111010;
      patterns[1313] = 50'b01_1110000110111111_1001111111111011_0100000111000100;
      patterns[1314] = 50'b10_1110000110111111_1001111111111011_1000000110111011;
      patterns[1315] = 50'b11_1110000110111111_1001111111111011_1111111111111111;
      patterns[1316] = 50'b00_1000010010100101_1111110001001000_1000000011101101;
      patterns[1317] = 50'b01_1000010010100101_1111110001001000_1000100001011101;
      patterns[1318] = 50'b10_1000010010100101_1111110001001000_1000010000000000;
      patterns[1319] = 50'b11_1000010010100101_1111110001001000_1111110011101101;
      patterns[1320] = 50'b00_0000101011000010_0001100000010110_0010001011011000;
      patterns[1321] = 50'b01_0000101011000010_0001100000010110_1111001010101100;
      patterns[1322] = 50'b10_0000101011000010_0001100000010110_0000100000000010;
      patterns[1323] = 50'b11_0000101011000010_0001100000010110_0001101011010110;
      patterns[1324] = 50'b00_0101111101010110_0011110000000000_1001101101010110;
      patterns[1325] = 50'b01_0101111101010110_0011110000000000_0010001101010110;
      patterns[1326] = 50'b10_0101111101010110_0011110000000000_0001110000000000;
      patterns[1327] = 50'b11_0101111101010110_0011110000000000_0111111101010110;
      patterns[1328] = 50'b00_1001000010010001_0000110001111111_1001110100010000;
      patterns[1329] = 50'b01_1001000010010001_0000110001111111_1000010000010010;
      patterns[1330] = 50'b10_1001000010010001_0000110001111111_0000000000010001;
      patterns[1331] = 50'b11_1001000010010001_0000110001111111_1001110011111111;
      patterns[1332] = 50'b00_1010000011001111_0000110011010110_1010110110100101;
      patterns[1333] = 50'b01_1010000011001111_0000110011010110_1001001111111001;
      patterns[1334] = 50'b10_1010000011001111_0000110011010110_0000000011000110;
      patterns[1335] = 50'b11_1010000011001111_0000110011010110_1010110011011111;
      patterns[1336] = 50'b00_0001011110011101_1101001100000101_1110101010100010;
      patterns[1337] = 50'b01_0001011110011101_1101001100000101_0100010010011000;
      patterns[1338] = 50'b10_0001011110011101_1101001100000101_0001001100000101;
      patterns[1339] = 50'b11_0001011110011101_1101001100000101_1101011110011101;
      patterns[1340] = 50'b00_1111011001001010_1010010011001011_1001101100010101;
      patterns[1341] = 50'b01_1111011001001010_1010010011001011_0101000101111111;
      patterns[1342] = 50'b10_1111011001001010_1010010011001011_1010010001001010;
      patterns[1343] = 50'b11_1111011001001010_1010010011001011_1111011011001011;
      patterns[1344] = 50'b00_1001000101100101_1000110011100101_0001111001001010;
      patterns[1345] = 50'b01_1001000101100101_1000110011100101_0000010010000000;
      patterns[1346] = 50'b10_1001000101100101_1000110011100101_1000000001100101;
      patterns[1347] = 50'b11_1001000101100101_1000110011100101_1001110111100101;
      patterns[1348] = 50'b00_1100010011111001_0101100110000010_0001111001111011;
      patterns[1349] = 50'b01_1100010011111001_0101100110000010_0110101101110111;
      patterns[1350] = 50'b10_1100010011111001_0101100110000010_0100000010000000;
      patterns[1351] = 50'b11_1100010011111001_0101100110000010_1101110111111011;
      patterns[1352] = 50'b00_0101100101101010_1101100011000010_0011001000101100;
      patterns[1353] = 50'b01_0101100101101010_1101100011000010_1000000010101000;
      patterns[1354] = 50'b10_0101100101101010_1101100011000010_0101100001000010;
      patterns[1355] = 50'b11_0101100101101010_1101100011000010_1101100111101010;
      patterns[1356] = 50'b00_1010010000010101_1011100011110010_0101110100000111;
      patterns[1357] = 50'b01_1010010000010101_1011100011110010_1110101100100011;
      patterns[1358] = 50'b10_1010010000010101_1011100011110010_1010000000010000;
      patterns[1359] = 50'b11_1010010000010101_1011100011110010_1011110011110111;
      patterns[1360] = 50'b00_0011011001100010_1100111111000001_0000011000100011;
      patterns[1361] = 50'b01_0011011001100010_1100111111000001_0110011010100001;
      patterns[1362] = 50'b10_0011011001100010_1100111111000001_0000011001000000;
      patterns[1363] = 50'b11_0011011001100010_1100111111000001_1111111111100011;
      patterns[1364] = 50'b00_0001100100100010_0000100010111100_0010000111011110;
      patterns[1365] = 50'b01_0001100100100010_0000100010111100_0001000001100110;
      patterns[1366] = 50'b10_0001100100100010_0000100010111100_0000100000100000;
      patterns[1367] = 50'b11_0001100100100010_0000100010111100_0001100110111110;
      patterns[1368] = 50'b00_1100010111101010_1001111110001001_0110010101110011;
      patterns[1369] = 50'b01_1100010111101010_1001111110001001_0010011001100001;
      patterns[1370] = 50'b10_1100010111101010_1001111110001001_1000010110001000;
      patterns[1371] = 50'b11_1100010111101010_1001111110001001_1101111111101011;
      patterns[1372] = 50'b00_0000011001010010_1001000010000110_1001011011011000;
      patterns[1373] = 50'b01_0000011001010010_1001000010000110_0111010111001100;
      patterns[1374] = 50'b10_0000011001010010_1001000010000110_0000000000000010;
      patterns[1375] = 50'b11_0000011001010010_1001000010000110_1001011011010110;
      patterns[1376] = 50'b00_1010011000110011_1100001001001110_0110100010000001;
      patterns[1377] = 50'b01_1010011000110011_1100001001001110_1110001111100101;
      patterns[1378] = 50'b10_1010011000110011_1100001001001110_1000001000000010;
      patterns[1379] = 50'b11_1010011000110011_1100001001001110_1110011001111111;
      patterns[1380] = 50'b00_1001110000001001_0111011100010011_0001001100011100;
      patterns[1381] = 50'b01_1001110000001001_0111011100010011_0010010011110110;
      patterns[1382] = 50'b10_1001110000001001_0111011100010011_0001010000000001;
      patterns[1383] = 50'b11_1001110000001001_0111011100010011_1111111100011011;
      patterns[1384] = 50'b00_1110011001011101_0010110100001100_0001001101101001;
      patterns[1385] = 50'b01_1110011001011101_0010110100001100_1011100101010001;
      patterns[1386] = 50'b10_1110011001011101_0010110100001100_0010010000001100;
      patterns[1387] = 50'b11_1110011001011101_0010110100001100_1110111101011101;
      patterns[1388] = 50'b00_1110011111101111_1000010011110111_0110110011100110;
      patterns[1389] = 50'b01_1110011111101111_1000010011110111_0110001011111000;
      patterns[1390] = 50'b10_1110011111101111_1000010011110111_1000010011100111;
      patterns[1391] = 50'b11_1110011111101111_1000010011110111_1110011111111111;
      patterns[1392] = 50'b00_1110001110000111_1100101110011100_1010111100100011;
      patterns[1393] = 50'b01_1110001110000111_1100101110011100_0001011111101011;
      patterns[1394] = 50'b10_1110001110000111_1100101110011100_1100001110000100;
      patterns[1395] = 50'b11_1110001110000111_1100101110011100_1110101110011111;
      patterns[1396] = 50'b00_0100110100100011_1101001100010111_0010000000111010;
      patterns[1397] = 50'b01_0100110100100011_1101001100010111_0111101000001100;
      patterns[1398] = 50'b10_0100110100100011_1101001100010111_0100000100000011;
      patterns[1399] = 50'b11_0100110100100011_1101001100010111_1101111100110111;
      patterns[1400] = 50'b00_1011110110110110_0100100101011100_0000011100010010;
      patterns[1401] = 50'b01_1011110110110110_0100100101011100_0111010001011010;
      patterns[1402] = 50'b10_1011110110110110_0100100101011100_0000100100010100;
      patterns[1403] = 50'b11_1011110110110110_0100100101011100_1111110111111110;
      patterns[1404] = 50'b00_0100101001100110_0100011001011001_1001000010111111;
      patterns[1405] = 50'b01_0100101001100110_0100011001011001_0000010000001101;
      patterns[1406] = 50'b10_0100101001100110_0100011001011001_0100001001000000;
      patterns[1407] = 50'b11_0100101001100110_0100011001011001_0100111001111111;
      patterns[1408] = 50'b00_1111110100101111_0111010001110100_0111000110100011;
      patterns[1409] = 50'b01_1111110100101111_0111010001110100_1000100010111011;
      patterns[1410] = 50'b10_1111110100101111_0111010001110100_0111010000100100;
      patterns[1411] = 50'b11_1111110100101111_0111010001110100_1111110101111111;
      patterns[1412] = 50'b00_1111010001100000_1011110100110111_1011000110010111;
      patterns[1413] = 50'b01_1111010001100000_1011110100110111_0011011100101001;
      patterns[1414] = 50'b10_1111010001100000_1011110100110111_1011010000100000;
      patterns[1415] = 50'b11_1111010001100000_1011110100110111_1111110101110111;
      patterns[1416] = 50'b00_1101010111011001_1000000100001011_0101011011100100;
      patterns[1417] = 50'b01_1101010111011001_1000000100001011_0101010011001110;
      patterns[1418] = 50'b10_1101010111011001_1000000100001011_1000000100001001;
      patterns[1419] = 50'b11_1101010111011001_1000000100001011_1101010111011011;
      patterns[1420] = 50'b00_0111001101001101_1111111100010011_0111001001100000;
      patterns[1421] = 50'b01_0111001101001101_1111111100010011_0111010000111010;
      patterns[1422] = 50'b10_0111001101001101_1111111100010011_0111001100000001;
      patterns[1423] = 50'b11_0111001101001101_1111111100010011_1111111101011111;
      patterns[1424] = 50'b00_1011001111000011_0001000011101111_1100010010110010;
      patterns[1425] = 50'b01_1011001111000011_0001000011101111_1010001011010100;
      patterns[1426] = 50'b10_1011001111000011_0001000011101111_0001000011000011;
      patterns[1427] = 50'b11_1011001111000011_0001000011101111_1011001111101111;
      patterns[1428] = 50'b00_1010010011000000_1101000010001001_0111010101001001;
      patterns[1429] = 50'b01_1010010011000000_1101000010001001_1101010000110111;
      patterns[1430] = 50'b10_1010010011000000_1101000010001001_1000000010000000;
      patterns[1431] = 50'b11_1010010011000000_1101000010001001_1111010011001001;
      patterns[1432] = 50'b00_0110000011110000_0010101101111010_1000110001101010;
      patterns[1433] = 50'b01_0110000011110000_0010101101111010_0011010101110110;
      patterns[1434] = 50'b10_0110000011110000_0010101101111010_0010000001110000;
      patterns[1435] = 50'b11_0110000011110000_0010101101111010_0110101111111010;
      patterns[1436] = 50'b00_1011101100111000_0000101100001001_1100011001000001;
      patterns[1437] = 50'b01_1011101100111000_0000101100001001_1011000000101111;
      patterns[1438] = 50'b10_1011101100111000_0000101100001001_0000101100001000;
      patterns[1439] = 50'b11_1011101100111000_0000101100001001_1011101100111001;
      patterns[1440] = 50'b00_0010000111101000_0100000011000101_0110001010101101;
      patterns[1441] = 50'b01_0010000111101000_0100000011000101_1110000100100011;
      patterns[1442] = 50'b10_0010000111101000_0100000011000101_0000000011000000;
      patterns[1443] = 50'b11_0010000111101000_0100000011000101_0110000111101101;
      patterns[1444] = 50'b00_0101011011000100_0011100110001111_1001000001010011;
      patterns[1445] = 50'b01_0101011011000100_0011100110001111_0001110100110101;
      patterns[1446] = 50'b10_0101011011000100_0011100110001111_0001000010000100;
      patterns[1447] = 50'b11_0101011011000100_0011100110001111_0111111111001111;
      patterns[1448] = 50'b00_1001101111011000_1110101001100100_1000011000111100;
      patterns[1449] = 50'b01_1001101111011000_1110101001100100_1011000101110100;
      patterns[1450] = 50'b10_1001101111011000_1110101001100100_1000101001000000;
      patterns[1451] = 50'b11_1001101111011000_1110101001100100_1111101111111100;
      patterns[1452] = 50'b00_0001101011110000_0000011100110101_0010001000100101;
      patterns[1453] = 50'b01_0001101011110000_0000011100110101_0001001110111011;
      patterns[1454] = 50'b10_0001101011110000_0000011100110101_0000001000110000;
      patterns[1455] = 50'b11_0001101011110000_0000011100110101_0001111111110101;
      patterns[1456] = 50'b00_0011010000100000_0101101101001100_1000111101101100;
      patterns[1457] = 50'b01_0011010000100000_0101101101001100_1101100011010100;
      patterns[1458] = 50'b10_0011010000100000_0101101101001100_0001000000000000;
      patterns[1459] = 50'b11_0011010000100000_0101101101001100_0111111101101100;
      patterns[1460] = 50'b00_0011011110101101_1011111111101100_1111011110011001;
      patterns[1461] = 50'b01_0011011110101101_1011111111101100_0111011111000001;
      patterns[1462] = 50'b10_0011011110101101_1011111111101100_0011011110101100;
      patterns[1463] = 50'b11_0011011110101101_1011111111101100_1011111111101101;
      patterns[1464] = 50'b00_1101111010011111_0101011110010100_0011011000110011;
      patterns[1465] = 50'b01_1101111010011111_0101011110010100_1000011100001011;
      patterns[1466] = 50'b10_1101111010011111_0101011110010100_0101011010010100;
      patterns[1467] = 50'b11_1101111010011111_0101011110010100_1101111110011111;
      patterns[1468] = 50'b00_1011001111111111_0011111010110111_1111001010110110;
      patterns[1469] = 50'b01_1011001111111111_0011111010110111_0111010101001000;
      patterns[1470] = 50'b10_1011001111111111_0011111010110111_0011001010110111;
      patterns[1471] = 50'b11_1011001111111111_0011111010110111_1011111111111111;
      patterns[1472] = 50'b00_1111110100110001_0001110000101101_0001100101011110;
      patterns[1473] = 50'b01_1111110100110001_0001110000101101_1110000100000100;
      patterns[1474] = 50'b10_1111110100110001_0001110000101101_0001110000100001;
      patterns[1475] = 50'b11_1111110100110001_0001110000101101_1111110100111101;
      patterns[1476] = 50'b00_1000101010010000_1110100000001101_0111001010011101;
      patterns[1477] = 50'b01_1000101010010000_1110100000001101_1010001010000011;
      patterns[1478] = 50'b10_1000101010010000_1110100000001101_1000100000000000;
      patterns[1479] = 50'b11_1000101010010000_1110100000001101_1110101010011101;
      patterns[1480] = 50'b00_0000100000010010_1101010111010101_1101110111100111;
      patterns[1481] = 50'b01_0000100000010010_1101010111010101_0011001000111101;
      patterns[1482] = 50'b10_0000100000010010_1101010111010101_0000000000010000;
      patterns[1483] = 50'b11_0000100000010010_1101010111010101_1101110111010111;
      patterns[1484] = 50'b00_1101000110001011_1011101001011011_1000101111100110;
      patterns[1485] = 50'b01_1101000110001011_1011101001011011_0001011100110000;
      patterns[1486] = 50'b10_1101000110001011_1011101001011011_1001000000001011;
      patterns[1487] = 50'b11_1101000110001011_1011101001011011_1111101111011011;
      patterns[1488] = 50'b00_0011010000100110_0010010111001011_0101100111110001;
      patterns[1489] = 50'b01_0011010000100110_0010010111001011_0000111001011011;
      patterns[1490] = 50'b10_0011010000100110_0010010111001011_0010010000000010;
      patterns[1491] = 50'b11_0011010000100110_0010010111001011_0011010111101111;
      patterns[1492] = 50'b00_0011100001000000_0001000111000011_0100101000000011;
      patterns[1493] = 50'b01_0011100001000000_0001000111000011_0010011001111101;
      patterns[1494] = 50'b10_0011100001000000_0001000111000011_0001000001000000;
      patterns[1495] = 50'b11_0011100001000000_0001000111000011_0011100111000011;
      patterns[1496] = 50'b00_0011000101100101_1011101000010101_1110101101111010;
      patterns[1497] = 50'b01_0011000101100101_1011101000010101_0111011101010000;
      patterns[1498] = 50'b10_0011000101100101_1011101000010101_0011000000000101;
      patterns[1499] = 50'b11_0011000101100101_1011101000010101_1011101101110101;
      patterns[1500] = 50'b00_0001111010001110_0111011110001011_1001011000011001;
      patterns[1501] = 50'b01_0001111010001110_0111011110001011_1010011100000011;
      patterns[1502] = 50'b10_0001111010001110_0111011110001011_0001011010001010;
      patterns[1503] = 50'b11_0001111010001110_0111011110001011_0111111110001111;
      patterns[1504] = 50'b00_0110100011011000_0010111001011110_1001011100110110;
      patterns[1505] = 50'b01_0110100011011000_0010111001011110_0011101001111010;
      patterns[1506] = 50'b10_0110100011011000_0010111001011110_0010100001011000;
      patterns[1507] = 50'b11_0110100011011000_0010111001011110_0110111011011110;
      patterns[1508] = 50'b00_0110101100001011_1011100011011011_0010001111100110;
      patterns[1509] = 50'b01_0110101100001011_1011100011011011_1011001000110000;
      patterns[1510] = 50'b10_0110101100001011_1011100011011011_0010100000001011;
      patterns[1511] = 50'b11_0110101100001011_1011100011011011_1111101111011011;
      patterns[1512] = 50'b00_1101011011101101_0100000110111001_0001100010100110;
      patterns[1513] = 50'b01_1101011011101101_0100000110111001_1001010100110100;
      patterns[1514] = 50'b10_1101011011101101_0100000110111001_0100000010101001;
      patterns[1515] = 50'b11_1101011011101101_0100000110111001_1101011111111101;
      patterns[1516] = 50'b00_0000111001011011_1000101111000001_1001101000011100;
      patterns[1517] = 50'b01_0000111001011011_1000101111000001_1000001010011010;
      patterns[1518] = 50'b10_0000111001011011_1000101111000001_0000101001000001;
      patterns[1519] = 50'b11_0000111001011011_1000101111000001_1000111111011011;
      patterns[1520] = 50'b00_1011110000010111_1110110011001010_1010100011100001;
      patterns[1521] = 50'b01_1011110000010111_1110110011001010_1100111101001101;
      patterns[1522] = 50'b10_1011110000010111_1110110011001010_1010110000000010;
      patterns[1523] = 50'b11_1011110000010111_1110110011001010_1111110011011111;
      patterns[1524] = 50'b00_1101001101001001_0011110010011100_0000111111100101;
      patterns[1525] = 50'b01_1101001101001001_0011110010011100_1001011010101101;
      patterns[1526] = 50'b10_1101001101001001_0011110010011100_0001000000001000;
      patterns[1527] = 50'b11_1101001101001001_0011110010011100_1111111111011101;
      patterns[1528] = 50'b00_1110001011101111_0000101100101101_1110111000011100;
      patterns[1529] = 50'b01_1110001011101111_0000101100101101_1101011111000010;
      patterns[1530] = 50'b10_1110001011101111_0000101100101101_0000001000101101;
      patterns[1531] = 50'b11_1110001011101111_0000101100101101_1110101111101111;
      patterns[1532] = 50'b00_1011010001110110_0011100101011111_1110110111010101;
      patterns[1533] = 50'b01_1011010001110110_0011100101011111_0111101100010111;
      patterns[1534] = 50'b10_1011010001110110_0011100101011111_0011000001010110;
      patterns[1535] = 50'b11_1011010001110110_0011100101011111_1011110101111111;
      patterns[1536] = 50'b00_0010100001011111_0001101000011011_0100001001111010;
      patterns[1537] = 50'b01_0010100001011111_0001101000011011_0000111001000100;
      patterns[1538] = 50'b10_0010100001011111_0001101000011011_0000100000011011;
      patterns[1539] = 50'b11_0010100001011111_0001101000011011_0011101001011111;
      patterns[1540] = 50'b00_0111000111000011_1101001101001000_0100010100001011;
      patterns[1541] = 50'b01_0111000111000011_1101001101001000_1001111001111011;
      patterns[1542] = 50'b10_0111000111000011_1101001101001000_0101000101000000;
      patterns[1543] = 50'b11_0111000111000011_1101001101001000_1111001111001011;
      patterns[1544] = 50'b00_0100011101111111_0000010110011010_0100110100011001;
      patterns[1545] = 50'b01_0100011101111111_0000010110011010_0100000111100101;
      patterns[1546] = 50'b10_0100011101111111_0000010110011010_0000010100011010;
      patterns[1547] = 50'b11_0100011101111111_0000010110011010_0100011111111111;
      patterns[1548] = 50'b00_1000100011000110_0011101100001001_1100001111001111;
      patterns[1549] = 50'b01_1000100011000110_0011101100001001_0100110110111101;
      patterns[1550] = 50'b10_1000100011000110_0011101100001001_0000100000000000;
      patterns[1551] = 50'b11_1000100011000110_0011101100001001_1011101111001111;
      patterns[1552] = 50'b00_1010100000101000_0001110011000010_1100010011101010;
      patterns[1553] = 50'b01_1010100000101000_0001110011000010_1000101101100110;
      patterns[1554] = 50'b10_1010100000101000_0001110011000010_0000100000000000;
      patterns[1555] = 50'b11_1010100000101000_0001110011000010_1011110011101010;
      patterns[1556] = 50'b00_0000010011101100_1000111010000000_1001001101101100;
      patterns[1557] = 50'b01_0000010011101100_1000111010000000_0111011001101100;
      patterns[1558] = 50'b10_0000010011101100_1000111010000000_0000010010000000;
      patterns[1559] = 50'b11_0000010011101100_1000111010000000_1000111011101100;
      patterns[1560] = 50'b00_0001010001111000_0000110011011111_0010000101010111;
      patterns[1561] = 50'b01_0001010001111000_0000110011011111_0000011110011001;
      patterns[1562] = 50'b10_0001010001111000_0000110011011111_0000010001011000;
      patterns[1563] = 50'b11_0001010001111000_0000110011011111_0001110011111111;
      patterns[1564] = 50'b00_1101010100011000_1100101001101000_1001111110000000;
      patterns[1565] = 50'b01_1101010100011000_1100101001101000_0000101010110000;
      patterns[1566] = 50'b10_1101010100011000_1100101001101000_1100000000001000;
      patterns[1567] = 50'b11_1101010100011000_1100101001101000_1101111101111000;
      patterns[1568] = 50'b00_1100011010111101_0011001010000000_1111100100111101;
      patterns[1569] = 50'b01_1100011010111101_0011001010000000_1001010000111101;
      patterns[1570] = 50'b10_1100011010111101_0011001010000000_0000001010000000;
      patterns[1571] = 50'b11_1100011010111101_0011001010000000_1111011010111101;
      patterns[1572] = 50'b00_0111010111101010_1001010110101111_0000101110011001;
      patterns[1573] = 50'b01_0111010111101010_1001010110101111_1110000000111011;
      patterns[1574] = 50'b10_0111010111101010_1001010110101111_0001010110101010;
      patterns[1575] = 50'b11_0111010111101010_1001010110101111_1111010111101111;
      patterns[1576] = 50'b00_0011011010000100_1010011010110100_1101110100111000;
      patterns[1577] = 50'b01_0011011010000100_1010011010110100_1000111111010000;
      patterns[1578] = 50'b10_0011011010000100_1010011010110100_0010011010000100;
      patterns[1579] = 50'b11_0011011010000100_1010011010110100_1011011010110100;
      patterns[1580] = 50'b00_1100100011110010_0010011101100110_1111000001011000;
      patterns[1581] = 50'b01_1100100011110010_0010011101100110_1010000110001100;
      patterns[1582] = 50'b10_1100100011110010_0010011101100110_0000000001100010;
      patterns[1583] = 50'b11_1100100011110010_0010011101100110_1110111111110110;
      patterns[1584] = 50'b00_0110100010111011_0010111000001000_1001011011000011;
      patterns[1585] = 50'b01_0110100010111011_0010111000001000_0011101010110011;
      patterns[1586] = 50'b10_0110100010111011_0010111000001000_0010100000001000;
      patterns[1587] = 50'b11_0110100010111011_0010111000001000_0110111010111011;
      patterns[1588] = 50'b00_1110001001111011_1111101101011001_1101110111010100;
      patterns[1589] = 50'b01_1110001001111011_1111101101011001_1110011100100010;
      patterns[1590] = 50'b10_1110001001111011_1111101101011001_1110001001011001;
      patterns[1591] = 50'b11_1110001001111011_1111101101011001_1111101101111011;
      patterns[1592] = 50'b00_0100110000111011_1001011000000110_1110001001000001;
      patterns[1593] = 50'b01_0100110000111011_1001011000000110_1011011000110101;
      patterns[1594] = 50'b10_0100110000111011_1001011000000110_0000010000000010;
      patterns[1595] = 50'b11_0100110000111011_1001011000000110_1101111000111111;
      patterns[1596] = 50'b00_0111000011000010_1010010011011111_0001010110100001;
      patterns[1597] = 50'b01_0111000011000010_1010010011011111_1100101111100011;
      patterns[1598] = 50'b10_0111000011000010_1010010011011111_0010000011000010;
      patterns[1599] = 50'b11_0111000011000010_1010010011011111_1111010011011111;
      patterns[1600] = 50'b00_1101100100010000_0001110101001111_1111011001011111;
      patterns[1601] = 50'b01_1101100100010000_0001110101001111_1011101111000001;
      patterns[1602] = 50'b10_1101100100010000_0001110101001111_0001100100000000;
      patterns[1603] = 50'b11_1101100100010000_0001110101001111_1101110101011111;
      patterns[1604] = 50'b00_0010000010101010_1101001001100110_1111001100010000;
      patterns[1605] = 50'b01_0010000010101010_1101001001100110_0100111001000100;
      patterns[1606] = 50'b10_0010000010101010_1101001001100110_0000000000100010;
      patterns[1607] = 50'b11_0010000010101010_1101001001100110_1111001011101110;
      patterns[1608] = 50'b00_0011111001010111_0011100110000100_0111011111011011;
      patterns[1609] = 50'b01_0011111001010111_0011100110000100_0000010011010011;
      patterns[1610] = 50'b10_0011111001010111_0011100110000100_0011100000000100;
      patterns[1611] = 50'b11_0011111001010111_0011100110000100_0011111111010111;
      patterns[1612] = 50'b00_0000110101011011_0111111111000011_1000110100011110;
      patterns[1613] = 50'b01_0000110101011011_0111111111000011_1000110110011000;
      patterns[1614] = 50'b10_0000110101011011_0111111111000011_0000110101000011;
      patterns[1615] = 50'b11_0000110101011011_0111111111000011_0111111111011011;
      patterns[1616] = 50'b00_0110011110011011_0110110110011011_1101010100110110;
      patterns[1617] = 50'b01_0110011110011011_0110110110011011_1111101000000000;
      patterns[1618] = 50'b10_0110011110011011_0110110110011011_0110010110011011;
      patterns[1619] = 50'b11_0110011110011011_0110110110011011_0110111110011011;
      patterns[1620] = 50'b00_1101100101010011_0110100001011111_0100000110110010;
      patterns[1621] = 50'b01_1101100101010011_0110100001011111_0111000011110100;
      patterns[1622] = 50'b10_1101100101010011_0110100001011111_0100100001010011;
      patterns[1623] = 50'b11_1101100101010011_0110100001011111_1111100101011111;
      patterns[1624] = 50'b00_1000011111110101_1110101001100001_0111001001010110;
      patterns[1625] = 50'b01_1000011111110101_1110101001100001_1001110110010100;
      patterns[1626] = 50'b10_1000011111110101_1110101001100001_1000001001100001;
      patterns[1627] = 50'b11_1000011111110101_1110101001100001_1110111111110101;
      patterns[1628] = 50'b00_1000100011001010_0000010110101110_1000111001111000;
      patterns[1629] = 50'b01_1000100011001010_0000010110101110_1000001100011100;
      patterns[1630] = 50'b10_1000100011001010_0000010110101110_0000000010001010;
      patterns[1631] = 50'b11_1000100011001010_0000010110101110_1000110111101110;
      patterns[1632] = 50'b00_0010011001011011_0110001000111000_1000100010010011;
      patterns[1633] = 50'b01_0010011001011011_0110001000111000_1100010000100011;
      patterns[1634] = 50'b10_0010011001011011_0110001000111000_0010001000011000;
      patterns[1635] = 50'b11_0010011001011011_0110001000111000_0110011001111011;
      patterns[1636] = 50'b00_1001011010000110_1100100110100001_0110000000100111;
      patterns[1637] = 50'b01_1001011010000110_1100100110100001_1100110011100101;
      patterns[1638] = 50'b10_1001011010000110_1100100110100001_1000000010000000;
      patterns[1639] = 50'b11_1001011010000110_1100100110100001_1101111110100111;
      patterns[1640] = 50'b00_0101101111110001_1101000001001110_0010110000111111;
      patterns[1641] = 50'b01_0101101111110001_1101000001001110_1000101110100011;
      patterns[1642] = 50'b10_0101101111110001_1101000001001110_0101000001000000;
      patterns[1643] = 50'b11_0101101111110001_1101000001001110_1101101111111111;
      patterns[1644] = 50'b00_0000010101110111_1100111111110010_1101010101101001;
      patterns[1645] = 50'b01_0000010101110111_1100111111110010_0011010110000101;
      patterns[1646] = 50'b10_0000010101110111_1100111111110010_0000010101110010;
      patterns[1647] = 50'b11_0000010101110111_1100111111110010_1100111111110111;
      patterns[1648] = 50'b00_1001001000110011_1111001011101110_1000010100100001;
      patterns[1649] = 50'b01_1001001000110011_1111001011101110_1001111101000101;
      patterns[1650] = 50'b10_1001001000110011_1111001011101110_1001001000100010;
      patterns[1651] = 50'b11_1001001000110011_1111001011101110_1111001011111111;
      patterns[1652] = 50'b00_0110001010110010_1111010010000000_0101011100110010;
      patterns[1653] = 50'b01_0110001010110010_1111010010000000_0110111000110010;
      patterns[1654] = 50'b10_0110001010110010_1111010010000000_0110000010000000;
      patterns[1655] = 50'b11_0110001010110010_1111010010000000_1111011010110010;
      patterns[1656] = 50'b00_0001010001010110_1101111110011110_1111001111110100;
      patterns[1657] = 50'b01_0001010001010110_1101111110011110_0011010010111000;
      patterns[1658] = 50'b10_0001010001010110_1101111110011110_0001010000010110;
      patterns[1659] = 50'b11_0001010001010110_1101111110011110_1101111111011110;
      patterns[1660] = 50'b00_1100010010100111_0001100000011000_1101110010111111;
      patterns[1661] = 50'b01_1100010010100111_0001100000011000_1010110010001111;
      patterns[1662] = 50'b10_1100010010100111_0001100000011000_0000000000000000;
      patterns[1663] = 50'b11_1100010010100111_0001100000011000_1101110010111111;
      patterns[1664] = 50'b00_0011010001000000_0110011100100010_1001101101100010;
      patterns[1665] = 50'b01_0011010001000000_0110011100100010_1100110100011110;
      patterns[1666] = 50'b10_0011010001000000_0110011100100010_0010010000000000;
      patterns[1667] = 50'b11_0011010001000000_0110011100100010_0111011101100010;
      patterns[1668] = 50'b00_1101010110101111_0110000001100010_0011011000010001;
      patterns[1669] = 50'b01_1101010110101111_0110000001100010_0111010101001101;
      patterns[1670] = 50'b10_1101010110101111_0110000001100010_0100000000100010;
      patterns[1671] = 50'b11_1101010110101111_0110000001100010_1111010111101111;
      patterns[1672] = 50'b00_1001100011011110_1111011010101010_1000111110001000;
      patterns[1673] = 50'b01_1001100011011110_1111011010101010_1010001000110100;
      patterns[1674] = 50'b10_1001100011011110_1111011010101010_1001000010001010;
      patterns[1675] = 50'b11_1001100011011110_1111011010101010_1111111011111110;
      patterns[1676] = 50'b00_1110000101000110_0110101011010001_0100110000010111;
      patterns[1677] = 50'b01_1110000101000110_0110101011010001_0111011001110101;
      patterns[1678] = 50'b10_1110000101000110_0110101011010001_0110000001000000;
      patterns[1679] = 50'b11_1110000101000110_0110101011010001_1110101111010111;
      patterns[1680] = 50'b00_1000100011001001_0100001010110001_1100101101111010;
      patterns[1681] = 50'b01_1000100011001001_0100001010110001_0100011000011000;
      patterns[1682] = 50'b10_1000100011001001_0100001010110001_0000000010000001;
      patterns[1683] = 50'b11_1000100011001001_0100001010110001_1100101011111001;
      patterns[1684] = 50'b00_1010110010010010_1011110111001011_0110101001011101;
      patterns[1685] = 50'b01_1010110010010010_1011110111001011_1110111011000111;
      patterns[1686] = 50'b10_1010110010010010_1011110111001011_1010110010000010;
      patterns[1687] = 50'b11_1010110010010010_1011110111001011_1011110111011011;
      patterns[1688] = 50'b00_1010100110000101_0100111101100001_1111100011100110;
      patterns[1689] = 50'b01_1010100110000101_0100111101100001_0101101000100100;
      patterns[1690] = 50'b10_1010100110000101_0100111101100001_0000100100000001;
      patterns[1691] = 50'b11_1010100110000101_0100111101100001_1110111111100101;
      patterns[1692] = 50'b00_1001110000001011_0011111001100010_1101101001101101;
      patterns[1693] = 50'b01_1001110000001011_0011111001100010_0101110110101001;
      patterns[1694] = 50'b10_1001110000001011_0011111001100010_0001110000000010;
      patterns[1695] = 50'b11_1001110000001011_0011111001100010_1011111001101011;
      patterns[1696] = 50'b00_1011100010111001_0101100101111010_0001001000110011;
      patterns[1697] = 50'b01_1011100010111001_0101100101111010_0101111100111111;
      patterns[1698] = 50'b10_1011100010111001_0101100101111010_0001100000111000;
      patterns[1699] = 50'b11_1011100010111001_0101100101111010_1111100111111011;
      patterns[1700] = 50'b00_0100100101011111_0001010001011111_0101110110111110;
      patterns[1701] = 50'b01_0100100101011111_0001010001011111_0011010100000000;
      patterns[1702] = 50'b10_0100100101011111_0001010001011111_0000000001011111;
      patterns[1703] = 50'b11_0100100101011111_0001010001011111_0101110101011111;
      patterns[1704] = 50'b00_0011101000111000_1011101000001110_1111010001000110;
      patterns[1705] = 50'b01_0011101000111000_1011101000001110_1000000000101010;
      patterns[1706] = 50'b10_0011101000111000_1011101000001110_0011101000001000;
      patterns[1707] = 50'b11_0011101000111000_1011101000001110_1011101000111110;
      patterns[1708] = 50'b00_0011010111110001_0011000101111000_0110011101101001;
      patterns[1709] = 50'b01_0011010111110001_0011000101111000_0000010001111001;
      patterns[1710] = 50'b10_0011010111110001_0011000101111000_0011000101110000;
      patterns[1711] = 50'b11_0011010111110001_0011000101111000_0011010111111001;
      patterns[1712] = 50'b00_1111001010111001_0001111010011101_0001000101010110;
      patterns[1713] = 50'b01_1111001010111001_0001111010011101_1101010000011100;
      patterns[1714] = 50'b10_1111001010111001_0001111010011101_0001001010011001;
      patterns[1715] = 50'b11_1111001010111001_0001111010011101_1111111010111101;
      patterns[1716] = 50'b00_1011011110000101_1010001111011001_0101101101011110;
      patterns[1717] = 50'b01_1011011110000101_1010001111011001_0001001110101100;
      patterns[1718] = 50'b10_1011011110000101_1010001111011001_1010001110000001;
      patterns[1719] = 50'b11_1011011110000101_1010001111011001_1011011111011101;
      patterns[1720] = 50'b00_0100110010010000_0101011001010010_1010001011100010;
      patterns[1721] = 50'b01_0100110010010000_0101011001010010_1111011000111110;
      patterns[1722] = 50'b10_0100110010010000_0101011001010010_0100010000010000;
      patterns[1723] = 50'b11_0100110010010000_0101011001010010_0101111011010010;
      patterns[1724] = 50'b00_1001010111111101_1111011101111110_1000110101111011;
      patterns[1725] = 50'b01_1001010111111101_1111011101111110_1001111001111111;
      patterns[1726] = 50'b10_1001010111111101_1111011101111110_1001010101111100;
      patterns[1727] = 50'b11_1001010111111101_1111011101111110_1111011111111111;
      patterns[1728] = 50'b00_0111000011010010_1000010001110101_1111010101000111;
      patterns[1729] = 50'b01_0111000011010010_1000010001110101_1110110001011101;
      patterns[1730] = 50'b10_0111000011010010_1000010001110101_0000000001010000;
      patterns[1731] = 50'b11_0111000011010010_1000010001110101_1111010011110111;
      patterns[1732] = 50'b00_0001001000110101_0010110011110000_0011111100100101;
      patterns[1733] = 50'b01_0001001000110101_0010110011110000_1110010101000101;
      patterns[1734] = 50'b10_0001001000110101_0010110011110000_0000000000110000;
      patterns[1735] = 50'b11_0001001000110101_0010110011110000_0011111011110101;
      patterns[1736] = 50'b00_1111010010100011_1011111101010101_1011001111111000;
      patterns[1737] = 50'b01_1111010010100011_1011111101010101_0011010101001110;
      patterns[1738] = 50'b10_1111010010100011_1011111101010101_1011010000000001;
      patterns[1739] = 50'b11_1111010010100011_1011111101010101_1111111111110111;
      patterns[1740] = 50'b00_0011011101100011_0011011101011111_0110111011000010;
      patterns[1741] = 50'b01_0011011101100011_0011011101011111_0000000000000100;
      patterns[1742] = 50'b10_0011011101100011_0011011101011111_0011011101000011;
      patterns[1743] = 50'b11_0011011101100011_0011011101011111_0011011101111111;
      patterns[1744] = 50'b00_0111011110101101_0000001000111010_0111100111100111;
      patterns[1745] = 50'b01_0111011110101101_0000001000111010_0111010101110011;
      patterns[1746] = 50'b10_0111011110101101_0000001000111010_0000001000101000;
      patterns[1747] = 50'b11_0111011110101101_0000001000111010_0111011110111111;
      patterns[1748] = 50'b00_0110100110001100_1000011100111001_1111000011000101;
      patterns[1749] = 50'b01_0110100110001100_1000011100111001_1110001001010011;
      patterns[1750] = 50'b10_0110100110001100_1000011100111001_0000000100001000;
      patterns[1751] = 50'b11_0110100110001100_1000011100111001_1110111110111101;
      patterns[1752] = 50'b00_0111010111101110_1110000000100100_0101011000010010;
      patterns[1753] = 50'b01_0111010111101110_1110000000100100_1001010111001010;
      patterns[1754] = 50'b10_0111010111101110_1110000000100100_0110000000100100;
      patterns[1755] = 50'b11_0111010111101110_1110000000100100_1111010111101110;
      patterns[1756] = 50'b00_0001110011110011_1110000110111000_1111111010101011;
      patterns[1757] = 50'b01_0001110011110011_1110000110111000_0011101100111011;
      patterns[1758] = 50'b10_0001110011110011_1110000110111000_0000000010110000;
      patterns[1759] = 50'b11_0001110011110011_1110000110111000_1111110111111011;
      patterns[1760] = 50'b00_1101110001100011_1001010001100001_0111000011000100;
      patterns[1761] = 50'b01_1101110001100011_1001010001100001_0100100000000010;
      patterns[1762] = 50'b10_1101110001100011_1001010001100001_1001010001100001;
      patterns[1763] = 50'b11_1101110001100011_1001010001100001_1101110001100011;
      patterns[1764] = 50'b00_1000001110001110_1010100011110101_0010110010000011;
      patterns[1765] = 50'b01_1000001110001110_1010100011110101_1101101010011001;
      patterns[1766] = 50'b10_1000001110001110_1010100011110101_1000000010000100;
      patterns[1767] = 50'b11_1000001110001110_1010100011110101_1010101111111111;
      patterns[1768] = 50'b00_1010010101000111_1110010101001011_1000101010010010;
      patterns[1769] = 50'b01_1010010101000111_1110010101001011_1011111111111100;
      patterns[1770] = 50'b10_1010010101000111_1110010101001011_1010010101000011;
      patterns[1771] = 50'b11_1010010101000111_1110010101001011_1110010101001111;
      patterns[1772] = 50'b00_1100011011100100_1100001110001011_1000101001101111;
      patterns[1773] = 50'b01_1100011011100100_1100001110001011_0000001101011001;
      patterns[1774] = 50'b10_1100011011100100_1100001110001011_1100001010000000;
      patterns[1775] = 50'b11_1100011011100100_1100001110001011_1100011111101111;
      patterns[1776] = 50'b00_1101110111011100_1100110010101101_1010101010001001;
      patterns[1777] = 50'b01_1101110111011100_1100110010101101_0001000100101111;
      patterns[1778] = 50'b10_1101110111011100_1100110010101101_1100110010001100;
      patterns[1779] = 50'b11_1101110111011100_1100110010101101_1101110111111101;
      patterns[1780] = 50'b00_0001010111110101_1000010111011000_1001101111001101;
      patterns[1781] = 50'b01_0001010111110101_1000010111011000_1001000000011101;
      patterns[1782] = 50'b10_0001010111110101_1000010111011000_0000010111010000;
      patterns[1783] = 50'b11_0001010111110101_1000010111011000_1001010111111101;
      patterns[1784] = 50'b00_1111110011110101_0000000010011111_1111110110010100;
      patterns[1785] = 50'b01_1111110011110101_0000000010011111_1111110001010110;
      patterns[1786] = 50'b10_1111110011110101_0000000010011111_0000000010010101;
      patterns[1787] = 50'b11_1111110011110101_0000000010011111_1111110011111111;
      patterns[1788] = 50'b00_0110011111101101_0101101001011010_1100001001000111;
      patterns[1789] = 50'b01_0110011111101101_0101101001011010_0000110110010011;
      patterns[1790] = 50'b10_0110011111101101_0101101001011010_0100001001001000;
      patterns[1791] = 50'b11_0110011111101101_0101101001011010_0111111111111111;
      patterns[1792] = 50'b00_0101111011001011_0100011011101110_1010010110111001;
      patterns[1793] = 50'b01_0101111011001011_0100011011101110_0001011111011101;
      patterns[1794] = 50'b10_0101111011001011_0100011011101110_0100011011001010;
      patterns[1795] = 50'b11_0101111011001011_0100011011101110_0101111011101111;
      patterns[1796] = 50'b00_0101010111011011_0110100111000010_1011111110011101;
      patterns[1797] = 50'b01_0101010111011011_0110100111000010_1110110000011001;
      patterns[1798] = 50'b10_0101010111011011_0110100111000010_0100000111000010;
      patterns[1799] = 50'b11_0101010111011011_0110100111000010_0111110111011011;
      patterns[1800] = 50'b00_0000111111000111_1111010000111010_0000010000000001;
      patterns[1801] = 50'b01_0000111111000111_1111010000111010_0001101110001101;
      patterns[1802] = 50'b10_0000111111000111_1111010000111010_0000010000000010;
      patterns[1803] = 50'b11_0000111111000111_1111010000111010_1111111111111111;
      patterns[1804] = 50'b00_1101011010110010_0010111010111001_0000010101101011;
      patterns[1805] = 50'b01_1101011010110010_0010111010111001_1010011111111001;
      patterns[1806] = 50'b10_1101011010110010_0010111010111001_0000011010110000;
      patterns[1807] = 50'b11_1101011010110010_0010111010111001_1111111010111011;
      patterns[1808] = 50'b00_1100110100111011_0001011101111111_1110010010111010;
      patterns[1809] = 50'b01_1100110100111011_0001011101111111_1011010110111100;
      patterns[1810] = 50'b10_1100110100111011_0001011101111111_0000010100111011;
      patterns[1811] = 50'b11_1100110100111011_0001011101111111_1101111101111111;
      patterns[1812] = 50'b00_1111101000101111_1011010001101100_1010111010011011;
      patterns[1813] = 50'b01_1111101000101111_1011010001101100_0100010111000011;
      patterns[1814] = 50'b10_1111101000101111_1011010001101100_1011000000101100;
      patterns[1815] = 50'b11_1111101000101111_1011010001101100_1111111001101111;
      patterns[1816] = 50'b00_0100100001010100_1001100110101110_1110001000000010;
      patterns[1817] = 50'b01_0100100001010100_1001100110101110_1010111010100110;
      patterns[1818] = 50'b10_0100100001010100_1001100110101110_0000100000000100;
      patterns[1819] = 50'b11_0100100001010100_1001100110101110_1101100111111110;
      patterns[1820] = 50'b00_1111100010001011_0011101001011010_0011001011100101;
      patterns[1821] = 50'b01_1111100010001011_0011101001011010_1011111000110001;
      patterns[1822] = 50'b10_1111100010001011_0011101001011010_0011100000001010;
      patterns[1823] = 50'b11_1111100010001011_0011101001011010_1111101011011011;
      patterns[1824] = 50'b00_0100010010101010_0000100001110010_0100110100011100;
      patterns[1825] = 50'b01_0100010010101010_0000100001110010_0011110000111000;
      patterns[1826] = 50'b10_0100010010101010_0000100001110010_0000000000100010;
      patterns[1827] = 50'b11_0100010010101010_0000100001110010_0100110011111010;
      patterns[1828] = 50'b00_0000111000000011_0001101100001001_0010100100001100;
      patterns[1829] = 50'b01_0000111000000011_0001101100001001_1111001011111010;
      patterns[1830] = 50'b10_0000111000000011_0001101100001001_0000101000000001;
      patterns[1831] = 50'b11_0000111000000011_0001101100001001_0001111100001011;
      patterns[1832] = 50'b00_0010000100111101_1101101001101101_1111101110101010;
      patterns[1833] = 50'b01_0010000100111101_1101101001101101_0100011011010000;
      patterns[1834] = 50'b10_0010000100111101_1101101001101101_0000000000101101;
      patterns[1835] = 50'b11_0010000100111101_1101101001101101_1111101101111101;
      patterns[1836] = 50'b00_1010001010011001_0001111010000100_1100000100011101;
      patterns[1837] = 50'b01_1010001010011001_0001111010000100_1000010000010101;
      patterns[1838] = 50'b10_1010001010011001_0001111010000100_0000001010000000;
      patterns[1839] = 50'b11_1010001010011001_0001111010000100_1011111010011101;
      patterns[1840] = 50'b00_1011011111000001_1011101001101100_0111001000101101;
      patterns[1841] = 50'b01_1011011111000001_1011101001101100_1111110101010101;
      patterns[1842] = 50'b10_1011011111000001_1011101001101100_1011001001000000;
      patterns[1843] = 50'b11_1011011111000001_1011101001101100_1011111111101101;
      patterns[1844] = 50'b00_0010111110101011_1101010011011101_0000010010001000;
      patterns[1845] = 50'b01_0010111110101011_1101010011011101_0101101011001110;
      patterns[1846] = 50'b10_0010111110101011_1101010011011101_0000010010001001;
      patterns[1847] = 50'b11_0010111110101011_1101010011011101_1111111111111111;
      patterns[1848] = 50'b00_0100001110001111_1100111001100010_0001000111110001;
      patterns[1849] = 50'b01_0100001110001111_1100111001100010_0111010100101101;
      patterns[1850] = 50'b10_0100001110001111_1100111001100010_0100001000000010;
      patterns[1851] = 50'b11_0100001110001111_1100111001100010_1100111111101111;
      patterns[1852] = 50'b00_0010111000101111_0011000000000101_0101111000110100;
      patterns[1853] = 50'b01_0010111000101111_0011000000000101_1111111000101010;
      patterns[1854] = 50'b10_0010111000101111_0011000000000101_0010000000000101;
      patterns[1855] = 50'b11_0010111000101111_0011000000000101_0011111000101111;
      patterns[1856] = 50'b00_0010111010011001_1111111000111100_0010110011010101;
      patterns[1857] = 50'b01_0010111010011001_1111111000111100_0011000001011101;
      patterns[1858] = 50'b10_0010111010011001_1111111000111100_0010111000011000;
      patterns[1859] = 50'b11_0010111010011001_1111111000111100_1111111010111101;
      patterns[1860] = 50'b00_0001100110110110_0101011111000011_0111000101111001;
      patterns[1861] = 50'b01_0001100110110110_0101011111000011_1100000111110011;
      patterns[1862] = 50'b10_0001100110110110_0101011111000011_0001000110000010;
      patterns[1863] = 50'b11_0001100110110110_0101011111000011_0101111111110111;
      patterns[1864] = 50'b00_0011100000110100_1111010111000000_0010110111110100;
      patterns[1865] = 50'b01_0011100000110100_1111010111000000_0100001001110100;
      patterns[1866] = 50'b10_0011100000110100_1111010111000000_0011000000000000;
      patterns[1867] = 50'b11_0011100000110100_1111010111000000_1111110111110100;
      patterns[1868] = 50'b00_0011110110010010_1001110110010011_1101101100100101;
      patterns[1869] = 50'b01_0011110110010010_1001110110010011_1001111111111111;
      patterns[1870] = 50'b10_0011110110010010_1001110110010011_0001110110010010;
      patterns[1871] = 50'b11_0011110110010010_1001110110010011_1011110110010011;
      patterns[1872] = 50'b00_0110011010011010_1111110000100100_0110001010111110;
      patterns[1873] = 50'b01_0110011010011010_1111110000100100_0110101001110110;
      patterns[1874] = 50'b10_0110011010011010_1111110000100100_0110010000000000;
      patterns[1875] = 50'b11_0110011010011010_1111110000100100_1111111010111110;
      patterns[1876] = 50'b00_1001001010110001_1000100110101111_0001110001100000;
      patterns[1877] = 50'b01_1001001010110001_1000100110101111_0000100100000010;
      patterns[1878] = 50'b10_1001001010110001_1000100110101111_1000000010100001;
      patterns[1879] = 50'b11_1001001010110001_1000100110101111_1001101110111111;
      patterns[1880] = 50'b00_1001100101110111_1100001100000100_0101110001111011;
      patterns[1881] = 50'b01_1001100101110111_1100001100000100_1101011001110011;
      patterns[1882] = 50'b10_1001100101110111_1100001100000100_1000000100000100;
      patterns[1883] = 50'b11_1001100101110111_1100001100000100_1101101101110111;
      patterns[1884] = 50'b00_0110111000001110_0011010110100101_1010001110110011;
      patterns[1885] = 50'b01_0110111000001110_0011010110100101_0011100001101001;
      patterns[1886] = 50'b10_0110111000001110_0011010110100101_0010010000000100;
      patterns[1887] = 50'b11_0110111000001110_0011010110100101_0111111110101111;
      patterns[1888] = 50'b00_0110000011100110_1111110111010110_0101111010111100;
      patterns[1889] = 50'b01_0110000011100110_1111110111010110_0110001100010000;
      patterns[1890] = 50'b10_0110000011100110_1111110111010110_0110000011000110;
      patterns[1891] = 50'b11_0110000011100110_1111110111010110_1111110111110110;
      patterns[1892] = 50'b00_0010000011001010_1000110000011100_1010110011100110;
      patterns[1893] = 50'b01_0010000011001010_1000110000011100_1001010010101110;
      patterns[1894] = 50'b10_0010000011001010_1000110000011100_0000000000001000;
      patterns[1895] = 50'b11_0010000011001010_1000110000011100_1010110011011110;
      patterns[1896] = 50'b00_1111000110100010_1110101000101001_1101101111001011;
      patterns[1897] = 50'b01_1111000110100010_1110101000101001_0000011101111001;
      patterns[1898] = 50'b10_1111000110100010_1110101000101001_1110000000100000;
      patterns[1899] = 50'b11_1111000110100010_1110101000101001_1111101110101011;
      patterns[1900] = 50'b00_1111010001011000_1001000010111111_1000010100010111;
      patterns[1901] = 50'b01_1111010001011000_1001000010111111_0110001110011001;
      patterns[1902] = 50'b10_1111010001011000_1001000010111111_1001000000011000;
      patterns[1903] = 50'b11_1111010001011000_1001000010111111_1111010011111111;
      patterns[1904] = 50'b00_1010110001100011_1111000000100000_1001110010000011;
      patterns[1905] = 50'b01_1010110001100011_1111000000100000_1011110001000011;
      patterns[1906] = 50'b10_1010110001100011_1111000000100000_1010000000100000;
      patterns[1907] = 50'b11_1010110001100011_1111000000100000_1111110001100011;
      patterns[1908] = 50'b00_0001111000111100_1000011001110000_1010010010101100;
      patterns[1909] = 50'b01_0001111000111100_1000011001110000_1001011111001100;
      patterns[1910] = 50'b10_0001111000111100_1000011001110000_0000011000110000;
      patterns[1911] = 50'b11_0001111000111100_1000011001110000_1001111001111100;
      patterns[1912] = 50'b00_1011001110100110_0010101000010110_1101110110111100;
      patterns[1913] = 50'b01_1011001110100110_0010101000010110_1000100110010000;
      patterns[1914] = 50'b10_1011001110100110_0010101000010110_0010001000000110;
      patterns[1915] = 50'b11_1011001110100110_0010101000010110_1011101110110110;
      patterns[1916] = 50'b00_0110000001001111_1010010100101110_0000010101111101;
      patterns[1917] = 50'b01_0110000001001111_1010010100101110_1011101100100001;
      patterns[1918] = 50'b10_0110000001001111_1010010100101110_0010000000001110;
      patterns[1919] = 50'b11_0110000001001111_1010010100101110_1110010101101111;
      patterns[1920] = 50'b00_0111100001001101_1111000101010101_0110100110100010;
      patterns[1921] = 50'b01_0111100001001101_1111000101010101_1000011011111000;
      patterns[1922] = 50'b10_0111100001001101_1111000101010101_0111000001000101;
      patterns[1923] = 50'b11_0111100001001101_1111000101010101_1111100101011101;
      patterns[1924] = 50'b00_0000101110010110_0001010001011010_0001111111110000;
      patterns[1925] = 50'b01_0000101110010110_0001010001011010_1111011100111100;
      patterns[1926] = 50'b10_0000101110010110_0001010001011010_0000000000010010;
      patterns[1927] = 50'b11_0000101110010110_0001010001011010_0001111111011110;
      patterns[1928] = 50'b00_1111101011100010_1000010100111101_1000000000011111;
      patterns[1929] = 50'b01_1111101011100010_1000010100111101_0111010110100101;
      patterns[1930] = 50'b10_1111101011100010_1000010100111101_1000000000100000;
      patterns[1931] = 50'b11_1111101011100010_1000010100111101_1111111111111111;
      patterns[1932] = 50'b00_0000010100000101_0000100101000000_0000111001000101;
      patterns[1933] = 50'b01_0000010100000101_0000100101000000_1111101111000101;
      patterns[1934] = 50'b10_0000010100000101_0000100101000000_0000000100000000;
      patterns[1935] = 50'b11_0000010100000101_0000100101000000_0000110101000101;
      patterns[1936] = 50'b00_1011110001100110_1000000101100011_0011110111001001;
      patterns[1937] = 50'b01_1011110001100110_1000000101100011_0011101100000011;
      patterns[1938] = 50'b10_1011110001100110_1000000101100011_1000000001100010;
      patterns[1939] = 50'b11_1011110001100110_1000000101100011_1011110101100111;
      patterns[1940] = 50'b00_0011110011010011_0011110100011011_0111100111101110;
      patterns[1941] = 50'b01_0011110011010011_0011110100011011_1111111110111000;
      patterns[1942] = 50'b10_0011110011010011_0011110100011011_0011110000010011;
      patterns[1943] = 50'b11_0011110011010011_0011110100011011_0011110111011011;
      patterns[1944] = 50'b00_1111111011110110_0001111001101000_0001110101011110;
      patterns[1945] = 50'b01_1111111011110110_0001111001101000_1110000010001110;
      patterns[1946] = 50'b10_1111111011110110_0001111001101000_0001111001100000;
      patterns[1947] = 50'b11_1111111011110110_0001111001101000_1111111011111110;
      patterns[1948] = 50'b00_1100001000100110_0110100011101000_0010101100001110;
      patterns[1949] = 50'b01_1100001000100110_0110100011101000_0101100100111110;
      patterns[1950] = 50'b10_1100001000100110_0110100011101000_0100000000100000;
      patterns[1951] = 50'b11_1100001000100110_0110100011101000_1110101011101110;
      patterns[1952] = 50'b00_0000001110110011_0010100010011111_0010110001010010;
      patterns[1953] = 50'b01_0000001110110011_0010100010011111_1101101100010100;
      patterns[1954] = 50'b10_0000001110110011_0010100010011111_0000000010010011;
      patterns[1955] = 50'b11_0000001110110011_0010100010011111_0010101110111111;
      patterns[1956] = 50'b00_0011111001000111_0001100011001010_0101011100010001;
      patterns[1957] = 50'b01_0011111001000111_0001100011001010_0010010101111101;
      patterns[1958] = 50'b10_0011111001000111_0001100011001010_0001100001000010;
      patterns[1959] = 50'b11_0011111001000111_0001100011001010_0011111011001111;
      patterns[1960] = 50'b00_0110100010101110_0010111011000011_1001011101110001;
      patterns[1961] = 50'b01_0110100010101110_0010111011000011_0011100111101011;
      patterns[1962] = 50'b10_0110100010101110_0010111011000011_0010100010000010;
      patterns[1963] = 50'b11_0110100010101110_0010111011000011_0110111011101111;
      patterns[1964] = 50'b00_0010101110101011_1111001111011000_0001111110000011;
      patterns[1965] = 50'b01_0010101110101011_1111001111011000_0011011111010011;
      patterns[1966] = 50'b10_0010101110101011_1111001111011000_0010001110001000;
      patterns[1967] = 50'b11_0010101110101011_1111001111011000_1111101111111011;
      patterns[1968] = 50'b00_1010011011010001_1010101001001000_0101000100011001;
      patterns[1969] = 50'b01_1010011011010001_1010101001001000_1111110010001001;
      patterns[1970] = 50'b10_1010011011010001_1010101001001000_1010001001000000;
      patterns[1971] = 50'b11_1010011011010001_1010101001001000_1010111011011001;
      patterns[1972] = 50'b00_1000111001100011_1000100010001000_0001011011101011;
      patterns[1973] = 50'b01_1000111001100011_1000100010001000_0000010111011011;
      patterns[1974] = 50'b10_1000111001100011_1000100010001000_1000100000000000;
      patterns[1975] = 50'b11_1000111001100011_1000100010001000_1000111011101011;
      patterns[1976] = 50'b00_1111010011111111_1100101000010110_1011111100010101;
      patterns[1977] = 50'b01_1111010011111111_1100101000010110_0010101011101001;
      patterns[1978] = 50'b10_1111010011111111_1100101000010110_1100000000010110;
      patterns[1979] = 50'b11_1111010011111111_1100101000010110_1111111011111111;
      patterns[1980] = 50'b00_0100110011101001_1100100100010110_0001010111111111;
      patterns[1981] = 50'b01_0100110011101001_1100100100010110_1000001111010011;
      patterns[1982] = 50'b10_0100110011101001_1100100100010110_0100100000000000;
      patterns[1983] = 50'b11_0100110011101001_1100100100010110_1100110111111111;
      patterns[1984] = 50'b00_1000001011011110_0001011110110111_1001101010010101;
      patterns[1985] = 50'b01_1000001011011110_0001011110110111_0110101100100111;
      patterns[1986] = 50'b10_1000001011011110_0001011110110111_0000001010010110;
      patterns[1987] = 50'b11_1000001011011110_0001011110110111_1001011111111111;
      patterns[1988] = 50'b00_1000100101000011_1010011010101001_0010111111101100;
      patterns[1989] = 50'b01_1000100101000011_1010011010101001_1110001010011010;
      patterns[1990] = 50'b10_1000100101000011_1010011010101001_1000000000000001;
      patterns[1991] = 50'b11_1000100101000011_1010011010101001_1010111111101011;
      patterns[1992] = 50'b00_0001001100011000_0110011000110101_0111100101001101;
      patterns[1993] = 50'b01_0001001100011000_0110011000110101_1010110011100011;
      patterns[1994] = 50'b10_0001001100011000_0110011000110101_0000001000010000;
      patterns[1995] = 50'b11_0001001100011000_0110011000110101_0111011100111101;
      patterns[1996] = 50'b00_1000001111101101_1010010011111010_0010100011100111;
      patterns[1997] = 50'b01_1000001111101101_1010010011111010_1101111011110011;
      patterns[1998] = 50'b10_1000001111101101_1010010011111010_1000000011101000;
      patterns[1999] = 50'b11_1000001111101101_1010010011111010_1010011111111111;
      patterns[2000] = 50'b00_0111100111110011_0101100101001011_1101001100111110;
      patterns[2001] = 50'b01_0111100111110011_0101100101001011_0010000010101000;
      patterns[2002] = 50'b10_0111100111110011_0101100101001011_0101100101000011;
      patterns[2003] = 50'b11_0111100111110011_0101100101001011_0111100111111011;
      patterns[2004] = 50'b00_1010001100011100_1101001111010010_0111011011101110;
      patterns[2005] = 50'b01_1010001100011100_1101001111010010_1100111101001010;
      patterns[2006] = 50'b10_1010001100011100_1101001111010010_1000001100010000;
      patterns[2007] = 50'b11_1010001100011100_1101001111010010_1111001111011110;
      patterns[2008] = 50'b00_0110101010001100_0101101010011101_1100010100101001;
      patterns[2009] = 50'b01_0110101010001100_0101101010011101_0000111111101111;
      patterns[2010] = 50'b10_0110101010001100_0101101010011101_0100101010001100;
      patterns[2011] = 50'b11_0110101010001100_0101101010011101_0111101010011101;
      patterns[2012] = 50'b00_0011001000110000_0101011010100110_1000100011010110;
      patterns[2013] = 50'b01_0011001000110000_0101011010100110_1101101110001010;
      patterns[2014] = 50'b10_0011001000110000_0101011010100110_0001001000100000;
      patterns[2015] = 50'b11_0011001000110000_0101011010100110_0111011010110110;
      patterns[2016] = 50'b00_0100101000110010_0000001000000101_0100110000110111;
      patterns[2017] = 50'b01_0100101000110010_0000001000000101_0100100000101101;
      patterns[2018] = 50'b10_0100101000110010_0000001000000101_0000001000000000;
      patterns[2019] = 50'b11_0100101000110010_0000001000000101_0100101000110111;
      patterns[2020] = 50'b00_0100111001111000_1000011000001100_1101010010000100;
      patterns[2021] = 50'b01_0100111001111000_1000011000001100_1100100001101100;
      patterns[2022] = 50'b10_0100111001111000_1000011000001100_0000011000001000;
      patterns[2023] = 50'b11_0100111001111000_1000011000001100_1100111001111100;
      patterns[2024] = 50'b00_0111011010000110_1100110101010000_0100001111010110;
      patterns[2025] = 50'b01_0111011010000110_1100110101010000_1010100100110110;
      patterns[2026] = 50'b10_0111011010000110_1100110101010000_0100010000000000;
      patterns[2027] = 50'b11_0111011010000110_1100110101010000_1111111111010110;
      patterns[2028] = 50'b00_0011111110011100_1100000111110011_0000000110001111;
      patterns[2029] = 50'b01_0011111110011100_1100000111110011_0111110110101001;
      patterns[2030] = 50'b10_0011111110011100_1100000111110011_0000000110010000;
      patterns[2031] = 50'b11_0011111110011100_1100000111110011_1111111111111111;
      patterns[2032] = 50'b00_1000100001110001_1000001011010110_0000101101000111;
      patterns[2033] = 50'b01_1000100001110001_1000001011010110_0000010110011011;
      patterns[2034] = 50'b10_1000100001110001_1000001011010110_1000000001010000;
      patterns[2035] = 50'b11_1000100001110001_1000001011010110_1000101011110111;
      patterns[2036] = 50'b00_0010101101000110_0011111011000101_0110101000001011;
      patterns[2037] = 50'b01_0010101101000110_0011111011000101_1110110010000001;
      patterns[2038] = 50'b10_0010101101000110_0011111011000101_0010101001000100;
      patterns[2039] = 50'b11_0010101101000110_0011111011000101_0011111111000111;
      patterns[2040] = 50'b00_1010001100011011_1100000111011100_0110010011110111;
      patterns[2041] = 50'b01_1010001100011011_1100000111011100_1110000100111111;
      patterns[2042] = 50'b10_1010001100011011_1100000111011100_1000000100011000;
      patterns[2043] = 50'b11_1010001100011011_1100000111011100_1110001111011111;
      patterns[2044] = 50'b00_1010110011101010_0111001011010010_0001111110111100;
      patterns[2045] = 50'b01_1010110011101010_0111001011010010_0011101000011000;
      patterns[2046] = 50'b10_1010110011101010_0111001011010010_0010000011000010;
      patterns[2047] = 50'b11_1010110011101010_0111001011010010_1111111011111010;
      patterns[2048] = 50'b00_1100101101101000_0001001010100101_1101111000001101;
      patterns[2049] = 50'b01_1100101101101000_0001001010100101_1011100011000011;
      patterns[2050] = 50'b10_1100101101101000_0001001010100101_0000001000100000;
      patterns[2051] = 50'b11_1100101101101000_0001001010100101_1101101111101101;
      patterns[2052] = 50'b00_0101101111000000_0100110011001101_1010100010001101;
      patterns[2053] = 50'b01_0101101111000000_0100110011001101_0000111011110011;
      patterns[2054] = 50'b10_0101101111000000_0100110011001101_0100100011000000;
      patterns[2055] = 50'b11_0101101111000000_0100110011001101_0101111111001101;
      patterns[2056] = 50'b00_1001100110101010_0011111110011011_1101100101000101;
      patterns[2057] = 50'b01_1001100110101010_0011111110011011_0101101000001111;
      patterns[2058] = 50'b10_1001100110101010_0011111110011011_0001100110001010;
      patterns[2059] = 50'b11_1001100110101010_0011111110011011_1011111110111011;
      patterns[2060] = 50'b00_1011001001001110_0000011100011011_1011100101101001;
      patterns[2061] = 50'b01_1011001001001110_0000011100011011_1010101100110011;
      patterns[2062] = 50'b10_1011001001001110_0000011100011011_0000001000001010;
      patterns[2063] = 50'b11_1011001001001110_0000011100011011_1011011101011111;
      patterns[2064] = 50'b00_0101010010000110_1110000000000110_0011010010001100;
      patterns[2065] = 50'b01_0101010010000110_1110000000000110_0111010010000000;
      patterns[2066] = 50'b10_0101010010000110_1110000000000110_0100000000000110;
      patterns[2067] = 50'b11_0101010010000110_1110000000000110_1111010010000110;
      patterns[2068] = 50'b00_0001110000100000_0011111101000011_0101101101100011;
      patterns[2069] = 50'b01_0001110000100000_0011111101000011_1101110011011101;
      patterns[2070] = 50'b10_0001110000100000_0011111101000011_0001110000000000;
      patterns[2071] = 50'b11_0001110000100000_0011111101000011_0011111101100011;
      patterns[2072] = 50'b00_1010100101010010_1100010000100100_0110110101110110;
      patterns[2073] = 50'b01_1010100101010010_1100010000100100_1110010100101110;
      patterns[2074] = 50'b10_1010100101010010_1100010000100100_1000000000000000;
      patterns[2075] = 50'b11_1010100101010010_1100010000100100_1110110101110110;
      patterns[2076] = 50'b00_0010011101111011_1111001111010101_0001101101010000;
      patterns[2077] = 50'b01_0010011101111011_1111001111010101_0011001110100110;
      patterns[2078] = 50'b10_0010011101111011_1111001111010101_0010001101010001;
      patterns[2079] = 50'b11_0010011101111011_1111001111010101_1111011111111111;
      patterns[2080] = 50'b00_1100001101001010_0110000110101010_0010010011110100;
      patterns[2081] = 50'b01_1100001101001010_0110000110101010_0110000110100000;
      patterns[2082] = 50'b10_1100001101001010_0110000110101010_0100000100001010;
      patterns[2083] = 50'b11_1100001101001010_0110000110101010_1110001111101010;
      patterns[2084] = 50'b00_1111101000110011_0010111001110100_0010100010100111;
      patterns[2085] = 50'b01_1111101000110011_0010111001110100_1100101110111111;
      patterns[2086] = 50'b10_1111101000110011_0010111001110100_0010101000110000;
      patterns[2087] = 50'b11_1111101000110011_0010111001110100_1111111001110111;
      patterns[2088] = 50'b00_0111100001111100_0111011011110011_1110111101101111;
      patterns[2089] = 50'b01_0111100001111100_0111011011110011_0000000110001001;
      patterns[2090] = 50'b10_0111100001111100_0111011011110011_0111000001110000;
      patterns[2091] = 50'b11_0111100001111100_0111011011110011_0111111011111111;
      patterns[2092] = 50'b00_0011000111111001_0110101011110101_1001110011101110;
      patterns[2093] = 50'b01_0011000111111001_0110101011110101_1100011100000100;
      patterns[2094] = 50'b10_0011000111111001_0110101011110101_0010000011110001;
      patterns[2095] = 50'b11_0011000111111001_0110101011110101_0111101111111101;
      patterns[2096] = 50'b00_1010000000111011_1101101001111000_0111101010110011;
      patterns[2097] = 50'b01_1010000000111011_1101101001111000_1100010111000011;
      patterns[2098] = 50'b10_1010000000111011_1101101001111000_1000000000111000;
      patterns[2099] = 50'b11_1010000000111011_1101101001111000_1111101001111011;
      patterns[2100] = 50'b00_0100100110110101_0011111110110011_1000100101101000;
      patterns[2101] = 50'b01_0100100110110101_0011111110110011_0000101000000010;
      patterns[2102] = 50'b10_0100100110110101_0011111110110011_0000100110110001;
      patterns[2103] = 50'b11_0100100110110101_0011111110110011_0111111110110111;
      patterns[2104] = 50'b00_0110110001111010_1101001101000001_0011111110111011;
      patterns[2105] = 50'b01_0110110001111010_1101001101000001_1001100100111001;
      patterns[2106] = 50'b10_0110110001111010_1101001101000001_0100000001000000;
      patterns[2107] = 50'b11_0110110001111010_1101001101000001_1111111101111011;
      patterns[2108] = 50'b00_0111011011010001_0110011010001010_1101110101011011;
      patterns[2109] = 50'b01_0111011011010001_0110011010001010_0001000001000111;
      patterns[2110] = 50'b10_0111011011010001_0110011010001010_0110011010000000;
      patterns[2111] = 50'b11_0111011011010001_0110011010001010_0111011011011011;
      patterns[2112] = 50'b00_1100110001101101_0110011001101100_0011001011011001;
      patterns[2113] = 50'b01_1100110001101101_0110011001101100_0110011000000001;
      patterns[2114] = 50'b10_1100110001101101_0110011001101100_0100010001101100;
      patterns[2115] = 50'b11_1100110001101101_0110011001101100_1110111001101101;
      patterns[2116] = 50'b00_1011001010000111_0000100100100000_1011101110100111;
      patterns[2117] = 50'b01_1011001010000111_0000100100100000_1010100101100111;
      patterns[2118] = 50'b10_1011001010000111_0000100100100000_0000000000000000;
      patterns[2119] = 50'b11_1011001010000111_0000100100100000_1011101110100111;
      patterns[2120] = 50'b00_0111010000110111_1011110100010011_0011000101001010;
      patterns[2121] = 50'b01_0111010000110111_1011110100010011_1011011100100100;
      patterns[2122] = 50'b10_0111010000110111_1011110100010011_0011010000010011;
      patterns[2123] = 50'b11_0111010000110111_1011110100010011_1111110100110111;
      patterns[2124] = 50'b00_0100110010001100_0001111001100010_0110101011101110;
      patterns[2125] = 50'b01_0100110010001100_0001111001100010_0010111000101010;
      patterns[2126] = 50'b10_0100110010001100_0001111001100010_0000110000000000;
      patterns[2127] = 50'b11_0100110010001100_0001111001100010_0101111011101110;
      patterns[2128] = 50'b00_0010001010011110_0010010100010011_0100011110110001;
      patterns[2129] = 50'b01_0010001010011110_0010010100010011_1111110110001011;
      patterns[2130] = 50'b10_0010001010011110_0010010100010011_0010000000010010;
      patterns[2131] = 50'b11_0010001010011110_0010010100010011_0010011110011111;
      patterns[2132] = 50'b00_1111010110111010_1011101001100111_1011000000100001;
      patterns[2133] = 50'b01_1111010110111010_1011101001100111_0011101101010011;
      patterns[2134] = 50'b10_1111010110111010_1011101001100111_1011000000100010;
      patterns[2135] = 50'b11_1111010110111010_1011101001100111_1111111111111111;
      patterns[2136] = 50'b00_0010001011111100_0011011001111111_0101100101111011;
      patterns[2137] = 50'b01_0010001011111100_0011011001111111_1110110001111101;
      patterns[2138] = 50'b10_0010001011111100_0011011001111111_0010001001111100;
      patterns[2139] = 50'b11_0010001011111100_0011011001111111_0011011011111111;
      patterns[2140] = 50'b00_1010101010000101_0110110100011111_0001011110100100;
      patterns[2141] = 50'b01_1010101010000101_0110110100011111_0011110101100110;
      patterns[2142] = 50'b10_1010101010000101_0110110100011111_0010100000000101;
      patterns[2143] = 50'b11_1010101010000101_0110110100011111_1110111110011111;
      patterns[2144] = 50'b00_1101011011101000_0101011011010011_0010110110111011;
      patterns[2145] = 50'b01_1101011011101000_0101011011010011_1000000000010101;
      patterns[2146] = 50'b10_1101011011101000_0101011011010011_0101011011000000;
      patterns[2147] = 50'b11_1101011011101000_0101011011010011_1101011011111011;
      patterns[2148] = 50'b00_0100011001100111_0010111101110001_0111010111011000;
      patterns[2149] = 50'b01_0100011001100111_0010111101110001_0001011011110110;
      patterns[2150] = 50'b10_0100011001100111_0010111101110001_0000011001100001;
      patterns[2151] = 50'b11_0100011001100111_0010111101110001_0110111101110111;
      patterns[2152] = 50'b00_0100100001001111_0010101000100000_0111001001101111;
      patterns[2153] = 50'b01_0100100001001111_0010101000100000_0001111000101111;
      patterns[2154] = 50'b10_0100100001001111_0010101000100000_0000100000000000;
      patterns[2155] = 50'b11_0100100001001111_0010101000100000_0110101001101111;
      patterns[2156] = 50'b00_1101001010001110_1110100111000101_1011110001010011;
      patterns[2157] = 50'b01_1101001010001110_1110100111000101_1110100011001001;
      patterns[2158] = 50'b10_1101001010001110_1110100111000101_1100000010000100;
      patterns[2159] = 50'b11_1101001010001110_1110100111000101_1111101111001111;
      patterns[2160] = 50'b00_0110001000000000_1000000111010001_1110001111010001;
      patterns[2161] = 50'b01_0110001000000000_1000000111010001_1110000000101111;
      patterns[2162] = 50'b10_0110001000000000_1000000111010001_0000000000000000;
      patterns[2163] = 50'b11_0110001000000000_1000000111010001_1110001111010001;
      patterns[2164] = 50'b00_1101001101100111_0101001000001001_0010010101110000;
      patterns[2165] = 50'b01_1101001101100111_0101001000001001_1000000101011110;
      patterns[2166] = 50'b10_1101001101100111_0101001000001001_0101001000000001;
      patterns[2167] = 50'b11_1101001101100111_0101001000001001_1101001101101111;
      patterns[2168] = 50'b00_0111000111011000_1111111110111101_0111000110010101;
      patterns[2169] = 50'b01_0111000111011000_1111111110111101_0111001000011011;
      patterns[2170] = 50'b10_0111000111011000_1111111110111101_0111000110011000;
      patterns[2171] = 50'b11_0111000111011000_1111111110111101_1111111111111101;
      patterns[2172] = 50'b00_1111000111101110_1011101010111000_1010110010100110;
      patterns[2173] = 50'b01_1111000111101110_1011101010111000_0011011100110110;
      patterns[2174] = 50'b10_1111000111101110_1011101010111000_1011000010101000;
      patterns[2175] = 50'b11_1111000111101110_1011101010111000_1111101111111110;
      patterns[2176] = 50'b00_0000010100010010_1111001110011110_1111100010110000;
      patterns[2177] = 50'b01_0000010100010010_1111001110011110_0001000101110100;
      patterns[2178] = 50'b10_0000010100010010_1111001110011110_0000000100010010;
      patterns[2179] = 50'b11_0000010100010010_1111001110011110_1111011110011110;
      patterns[2180] = 50'b00_0101111011001110_0110111101110101_1100111001000011;
      patterns[2181] = 50'b01_0101111011001110_0110111101110101_1110111101011001;
      patterns[2182] = 50'b10_0101111011001110_0110111101110101_0100111001000100;
      patterns[2183] = 50'b11_0101111011001110_0110111101110101_0111111111111111;
      patterns[2184] = 50'b00_0000010001101101_1111000000101111_1111010010011100;
      patterns[2185] = 50'b01_0000010001101101_1111000000101111_0001010000111110;
      patterns[2186] = 50'b10_0000010001101101_1111000000101111_0000000000101101;
      patterns[2187] = 50'b11_0000010001101101_1111000000101111_1111010001101111;
      patterns[2188] = 50'b00_0011011010101111_0110011100110000_1001110111011111;
      patterns[2189] = 50'b01_0011011010101111_0110011100110000_1100111101111111;
      patterns[2190] = 50'b10_0011011010101111_0110011100110000_0010011000100000;
      patterns[2191] = 50'b11_0011011010101111_0110011100110000_0111011110111111;
      patterns[2192] = 50'b00_0011001100101100_0011010010001001_0110011110110101;
      patterns[2193] = 50'b01_0011001100101100_0011010010001001_1111111010100011;
      patterns[2194] = 50'b10_0011001100101100_0011010010001001_0011000000001000;
      patterns[2195] = 50'b11_0011001100101100_0011010010001001_0011011110101101;
      patterns[2196] = 50'b00_0000000001001111_0110011100000011_0110011101010010;
      patterns[2197] = 50'b01_0000000001001111_0110011100000011_1001100101001100;
      patterns[2198] = 50'b10_0000000001001111_0110011100000011_0000000000000011;
      patterns[2199] = 50'b11_0000000001001111_0110011100000011_0110011101001111;
      patterns[2200] = 50'b00_1101100100011111_0100110101101110_0010011010001101;
      patterns[2201] = 50'b01_1101100100011111_0100110101101110_1000101110110001;
      patterns[2202] = 50'b10_1101100100011111_0100110101101110_0100100100001110;
      patterns[2203] = 50'b11_1101100100011111_0100110101101110_1101110101111111;
      patterns[2204] = 50'b00_0001011000111111_0010110000100000_0100001001011111;
      patterns[2205] = 50'b01_0001011000111111_0010110000100000_1110101000011111;
      patterns[2206] = 50'b10_0001011000111111_0010110000100000_0000010000100000;
      patterns[2207] = 50'b11_0001011000111111_0010110000100000_0011111000111111;
      patterns[2208] = 50'b00_0110110100111011_0100000110101111_1010111011101010;
      patterns[2209] = 50'b01_0110110100111011_0100000110101111_0010101110001100;
      patterns[2210] = 50'b10_0110110100111011_0100000110101111_0100000100101011;
      patterns[2211] = 50'b11_0110110100111011_0100000110101111_0110110110111111;
      patterns[2212] = 50'b00_0110111101011111_1101011010001101_0100010111101100;
      patterns[2213] = 50'b01_0110111101011111_1101011010001101_1001100011010010;
      patterns[2214] = 50'b10_0110111101011111_1101011010001101_0100011000001101;
      patterns[2215] = 50'b11_0110111101011111_1101011010001101_1111111111011111;
      patterns[2216] = 50'b00_1000101101101010_0011001111010111_1011111101000001;
      patterns[2217] = 50'b01_1000101101101010_0011001111010111_0101011110010011;
      patterns[2218] = 50'b10_1000101101101010_0011001111010111_0000001101000010;
      patterns[2219] = 50'b11_1000101101101010_0011001111010111_1011101111111111;
      patterns[2220] = 50'b00_1100001001101010_1001100110001111_0101101111111001;
      patterns[2221] = 50'b01_1100001001101010_1001100110001111_0010100011011011;
      patterns[2222] = 50'b10_1100001001101010_1001100110001111_1000000000001010;
      patterns[2223] = 50'b11_1100001001101010_1001100110001111_1101101111101111;
      patterns[2224] = 50'b00_0101110110100011_1010001010111010_0000000001011101;
      patterns[2225] = 50'b01_0101110110100011_1010001010111010_1011101011101001;
      patterns[2226] = 50'b10_0101110110100011_1010001010111010_0000000010100010;
      patterns[2227] = 50'b11_0101110110100011_1010001010111010_1111111110111011;
      patterns[2228] = 50'b00_0111001000111101_1010100111101010_0001110000100111;
      patterns[2229] = 50'b01_0111001000111101_1010100111101010_1100100001010011;
      patterns[2230] = 50'b10_0111001000111101_1010100111101010_0010000000101000;
      patterns[2231] = 50'b11_0111001000111101_1010100111101010_1111101111111111;
      patterns[2232] = 50'b00_1110010101101111_0101100110101001_0011111100011000;
      patterns[2233] = 50'b01_1110010101101111_0101100110101001_1000101111000110;
      patterns[2234] = 50'b10_1110010101101111_0101100110101001_0100000100101001;
      patterns[2235] = 50'b11_1110010101101111_0101100110101001_1111110111101111;
      patterns[2236] = 50'b00_0000100110100010_0111110101101011_1000011100001101;
      patterns[2237] = 50'b01_0000100110100010_0111110101101011_1000110000110111;
      patterns[2238] = 50'b10_0000100110100010_0111110101101011_0000100100100010;
      patterns[2239] = 50'b11_0000100110100010_0111110101101011_0111110111101011;
      patterns[2240] = 50'b00_0100000001100100_1011000001010101_1111000010111001;
      patterns[2241] = 50'b01_0100000001100100_1011000001010101_1001000000001111;
      patterns[2242] = 50'b10_0100000001100100_1011000001010101_0000000001000100;
      patterns[2243] = 50'b11_0100000001100100_1011000001010101_1111000001110101;
      patterns[2244] = 50'b00_0100111011000010_1011001001011011_0000000100011101;
      patterns[2245] = 50'b01_0100111011000010_1011001001011011_1001110001100111;
      patterns[2246] = 50'b10_0100111011000010_1011001001011011_0000001001000010;
      patterns[2247] = 50'b11_0100111011000010_1011001001011011_1111111011011011;
      patterns[2248] = 50'b00_0001011101000111_1111000110110001_0000100011111000;
      patterns[2249] = 50'b01_0001011101000111_1111000110110001_0010010110010110;
      patterns[2250] = 50'b10_0001011101000111_1111000110110001_0001000100000001;
      patterns[2251] = 50'b11_0001011101000111_1111000110110001_1111011111110111;
      patterns[2252] = 50'b00_0001111110011101_0110000011001100_1000000001101001;
      patterns[2253] = 50'b01_0001111110011101_0110000011001100_1011111011010001;
      patterns[2254] = 50'b10_0001111110011101_0110000011001100_0000000010001100;
      patterns[2255] = 50'b11_0001111110011101_0110000011001100_0111111111011101;
      patterns[2256] = 50'b00_1110010011010110_1010000001010101_1000010100101011;
      patterns[2257] = 50'b01_1110010011010110_1010000001010101_0100010010000001;
      patterns[2258] = 50'b10_1110010011010110_1010000001010101_1010000001010100;
      patterns[2259] = 50'b11_1110010011010110_1010000001010101_1110010011010111;
      patterns[2260] = 50'b00_0101101000001101_0010101011100111_1000010011110100;
      patterns[2261] = 50'b01_0101101000001101_0010101011100111_0010111100100110;
      patterns[2262] = 50'b10_0101101000001101_0010101011100111_0000101000000101;
      patterns[2263] = 50'b11_0101101000001101_0010101011100111_0111101011101111;
      patterns[2264] = 50'b00_1010011001101011_1101011000101111_0111110010011010;
      patterns[2265] = 50'b01_1010011001101011_1101011000101111_1101000000111100;
      patterns[2266] = 50'b10_1010011001101011_1101011000101111_1000011000101011;
      patterns[2267] = 50'b11_1010011001101011_1101011000101111_1111011001101111;
      patterns[2268] = 50'b00_0000101101001100_0001110010101000_0010011111110100;
      patterns[2269] = 50'b01_0000101101001100_0001110010101000_1110111010100100;
      patterns[2270] = 50'b10_0000101101001100_0001110010101000_0000100000001000;
      patterns[2271] = 50'b11_0000101101001100_0001110010101000_0001111111101100;
      patterns[2272] = 50'b00_1101010111111011_0010110010010100_0000001010001111;
      patterns[2273] = 50'b01_1101010111111011_0010110010010100_1010100101100111;
      patterns[2274] = 50'b10_1101010111111011_0010110010010100_0000010010010000;
      patterns[2275] = 50'b11_1101010111111011_0010110010010100_1111110111111111;
      patterns[2276] = 50'b00_0000001111111101_0100111010101100_0101001010101001;
      patterns[2277] = 50'b01_0000001111111101_0100111010101100_1011010101010001;
      patterns[2278] = 50'b10_0000001111111101_0100111010101100_0000001010101100;
      patterns[2279] = 50'b11_0000001111111101_0100111010101100_0100111111111101;
      patterns[2280] = 50'b00_0100001000101000_0111000011101010_1011001100010010;
      patterns[2281] = 50'b01_0100001000101000_0111000011101010_1101000100111110;
      patterns[2282] = 50'b10_0100001000101000_0111000011101010_0100000000101000;
      patterns[2283] = 50'b11_0100001000101000_0111000011101010_0111001011101010;
      patterns[2284] = 50'b00_1011011100011111_0100101100000001_0000001000100000;
      patterns[2285] = 50'b01_1011011100011111_0100101100000001_0110110000011110;
      patterns[2286] = 50'b10_1011011100011111_0100101100000001_0000001100000001;
      patterns[2287] = 50'b11_1011011100011111_0100101100000001_1111111100011111;
      patterns[2288] = 50'b00_0111011001011111_1110100110000101_0101111111100100;
      patterns[2289] = 50'b01_0111011001011111_1110100110000101_1000110011011010;
      patterns[2290] = 50'b10_0111011001011111_1110100110000101_0110000000000101;
      patterns[2291] = 50'b11_0111011001011111_1110100110000101_1111111111011111;
      patterns[2292] = 50'b00_1111101110000011_0110011000100011_0110000110100110;
      patterns[2293] = 50'b01_1111101110000011_0110011000100011_1001010101100000;
      patterns[2294] = 50'b10_1111101110000011_0110011000100011_0110001000000011;
      patterns[2295] = 50'b11_1111101110000011_0110011000100011_1111111110100011;
      patterns[2296] = 50'b00_1110101000110110_0001010101111010_1111111110110000;
      patterns[2297] = 50'b01_1110101000110110_0001010101111010_1101010010111100;
      patterns[2298] = 50'b10_1110101000110110_0001010101111010_0000000000110010;
      patterns[2299] = 50'b11_1110101000110110_0001010101111010_1111111101111110;
      patterns[2300] = 50'b00_1110000010011111_1001100110000101_0111101000100100;
      patterns[2301] = 50'b01_1110000010011111_1001100110000101_0100011100011010;
      patterns[2302] = 50'b10_1110000010011111_1001100110000101_1000000010000101;
      patterns[2303] = 50'b11_1110000010011111_1001100110000101_1111100110011111;
      patterns[2304] = 50'b00_0001110010010100_1010000101110011_1011111000000111;
      patterns[2305] = 50'b01_0001110010010100_1010000101110011_0111101100100001;
      patterns[2306] = 50'b10_0001110010010100_1010000101110011_0000000000010000;
      patterns[2307] = 50'b11_0001110010010100_1010000101110011_1011110111110111;
      patterns[2308] = 50'b00_0100100011001011_1111000001011110_0011100100101001;
      patterns[2309] = 50'b01_0100100011001011_1111000001011110_0101100001101101;
      patterns[2310] = 50'b10_0100100011001011_1111000001011110_0100000001001010;
      patterns[2311] = 50'b11_0100100011001011_1111000001011110_1111100011011111;
      patterns[2312] = 50'b00_0001010001001110_1100001011001001_1101011100010111;
      patterns[2313] = 50'b01_0001010001001110_1100001011001001_0101000110000101;
      patterns[2314] = 50'b10_0001010001001110_1100001011001001_0000000001001000;
      patterns[2315] = 50'b11_0001010001001110_1100001011001001_1101011011001111;
      patterns[2316] = 50'b00_0110010001011111_0100001010011101_1010011011111100;
      patterns[2317] = 50'b01_0110010001011111_0100001010011101_0010000111000010;
      patterns[2318] = 50'b10_0110010001011111_0100001010011101_0100000000011101;
      patterns[2319] = 50'b11_0110010001011111_0100001010011101_0110011011011111;
      patterns[2320] = 50'b00_0111110100111010_0100100101111100_1100011010110110;
      patterns[2321] = 50'b01_0111110100111010_0100100101111100_0011001110111110;
      patterns[2322] = 50'b10_0111110100111010_0100100101111100_0100100100111000;
      patterns[2323] = 50'b11_0111110100111010_0100100101111100_0111110101111110;
      patterns[2324] = 50'b00_0111101000101011_1100110100101111_0100011101011010;
      patterns[2325] = 50'b01_0111101000101011_1100110100101111_1010110011111100;
      patterns[2326] = 50'b10_0111101000101011_1100110100101111_0100100000101011;
      patterns[2327] = 50'b11_0111101000101011_1100110100101111_1111111100101111;
      patterns[2328] = 50'b00_1011110111101100_1000000011000010_0011111010101110;
      patterns[2329] = 50'b01_1011110111101100_1000000011000010_0011110100101010;
      patterns[2330] = 50'b10_1011110111101100_1000000011000010_1000000011000000;
      patterns[2331] = 50'b11_1011110111101100_1000000011000010_1011110111101110;
      patterns[2332] = 50'b00_1010001100111101_0011000111111011_1101010100111000;
      patterns[2333] = 50'b01_1010001100111101_0011000111111011_0111000101000010;
      patterns[2334] = 50'b10_1010001100111101_0011000111111011_0010000100111001;
      patterns[2335] = 50'b11_1010001100111101_0011000111111011_1011001111111111;
      patterns[2336] = 50'b00_1110111110100011_0110010101000000_0101010011100011;
      patterns[2337] = 50'b01_1110111110100011_0110010101000000_1000101001100011;
      patterns[2338] = 50'b10_1110111110100011_0110010101000000_0110010100000000;
      patterns[2339] = 50'b11_1110111110100011_0110010101000000_1110111111100011;
      patterns[2340] = 50'b00_0100000011111011_1000110101001110_1100111001001001;
      patterns[2341] = 50'b01_0100000011111011_1000110101001110_1011001110101101;
      patterns[2342] = 50'b10_0100000011111011_1000110101001110_0000000001001010;
      patterns[2343] = 50'b11_0100000011111011_1000110101001110_1100110111111111;
      patterns[2344] = 50'b00_1001011100010000_1100111100111010_0110011001001010;
      patterns[2345] = 50'b01_1001011100010000_1100111100111010_1100011111010110;
      patterns[2346] = 50'b10_1001011100010000_1100111100111010_1000011100010000;
      patterns[2347] = 50'b11_1001011100010000_1100111100111010_1101111100111010;
      patterns[2348] = 50'b00_1111110111111100_1001100110001111_1001011110001011;
      patterns[2349] = 50'b01_1111110111111100_1001100110001111_0110010001101101;
      patterns[2350] = 50'b10_1111110111111100_1001100110001111_1001100110001100;
      patterns[2351] = 50'b11_1111110111111100_1001100110001111_1111110111111111;
      patterns[2352] = 50'b00_0101101000000010_1110111000111011_0100100000111101;
      patterns[2353] = 50'b01_0101101000000010_1110111000111011_0110101111000111;
      patterns[2354] = 50'b10_0101101000000010_1110111000111011_0100101000000010;
      patterns[2355] = 50'b11_0101101000000010_1110111000111011_1111111000111011;
      patterns[2356] = 50'b00_0001101100101101_0100110101101110_0110100010011011;
      patterns[2357] = 50'b01_0001101100101101_0100110101101110_1100110110111111;
      patterns[2358] = 50'b10_0001101100101101_0100110101101110_0000100100101100;
      patterns[2359] = 50'b11_0001101100101101_0100110101101110_0101111101101111;
      patterns[2360] = 50'b00_1011001100100000_1101101100001001_1000111000101001;
      patterns[2361] = 50'b01_1011001100100000_1101101100001001_1101100000010111;
      patterns[2362] = 50'b10_1011001100100000_1101101100001001_1001001100000000;
      patterns[2363] = 50'b11_1011001100100000_1101101100001001_1111101100101001;
      patterns[2364] = 50'b00_1010010000101000_1111101111111010_1010000000100010;
      patterns[2365] = 50'b01_1010010000101000_1111101111111010_1010100000101110;
      patterns[2366] = 50'b10_1010010000101000_1111101111111010_1010000000101000;
      patterns[2367] = 50'b11_1010010000101000_1111101111111010_1111111111111010;
      patterns[2368] = 50'b00_1101001000111000_0001001111100000_1110011000011000;
      patterns[2369] = 50'b01_1101001000111000_0001001111100000_1011111001011000;
      patterns[2370] = 50'b10_1101001000111000_0001001111100000_0001001000100000;
      patterns[2371] = 50'b11_1101001000111000_0001001111100000_1101001111111000;
      patterns[2372] = 50'b00_1110011011000111_1100000101000010_1010100000001001;
      patterns[2373] = 50'b01_1110011011000111_1100000101000010_0010010110000101;
      patterns[2374] = 50'b10_1110011011000111_1100000101000010_1100000001000010;
      patterns[2375] = 50'b11_1110011011000111_1100000101000010_1110011111000111;
      patterns[2376] = 50'b00_0110110011010111_0110111001011000_1101101100101111;
      patterns[2377] = 50'b01_0110110011010111_0110111001011000_1111111001111111;
      patterns[2378] = 50'b10_0110110011010111_0110111001011000_0110110001010000;
      patterns[2379] = 50'b11_0110110011010111_0110111001011000_0110111011011111;
      patterns[2380] = 50'b00_0011001101011110_1111000101110000_0010010011001110;
      patterns[2381] = 50'b01_0011001101011110_1111000101110000_0100000111101110;
      patterns[2382] = 50'b10_0011001101011110_1111000101110000_0011000101010000;
      patterns[2383] = 50'b11_0011001101011110_1111000101110000_1111001101111110;
      patterns[2384] = 50'b00_0100000000101001_0110100101011100_1010100110000101;
      patterns[2385] = 50'b01_0100000000101001_0110100101011100_1101011011001101;
      patterns[2386] = 50'b10_0100000000101001_0110100101011100_0100000000001000;
      patterns[2387] = 50'b11_0100000000101001_0110100101011100_0110100101111101;
      patterns[2388] = 50'b00_0111110000101011_0101001110000000_1100111110101011;
      patterns[2389] = 50'b01_0111110000101011_0101001110000000_0010100010101011;
      patterns[2390] = 50'b10_0111110000101011_0101001110000000_0101000000000000;
      patterns[2391] = 50'b11_0111110000101011_0101001110000000_0111111110101011;
      patterns[2392] = 50'b00_0110101001001111_1101000100100100_0011101101110011;
      patterns[2393] = 50'b01_0110101001001111_1101000100100100_1001100100101011;
      patterns[2394] = 50'b10_0110101001001111_1101000100100100_0100000000000100;
      patterns[2395] = 50'b11_0110101001001111_1101000100100100_1111101101101111;
      patterns[2396] = 50'b00_1110001111011000_0010110000001111_0000111111100111;
      patterns[2397] = 50'b01_1110001111011000_0010110000001111_1011011111001001;
      patterns[2398] = 50'b10_1110001111011000_0010110000001111_0010000000001000;
      patterns[2399] = 50'b11_1110001111011000_0010110000001111_1110111111011111;
      patterns[2400] = 50'b00_1000111010110100_0101011000010110_1110010011001010;
      patterns[2401] = 50'b01_1000111010110100_0101011000010110_0011100010011110;
      patterns[2402] = 50'b10_1000111010110100_0101011000010110_0000011000010100;
      patterns[2403] = 50'b11_1000111010110100_0101011000010110_1101111010110110;
      patterns[2404] = 50'b00_1010110000110000_0111111111010000_0010110000000000;
      patterns[2405] = 50'b01_1010110000110000_0111111111010000_0010110001100000;
      patterns[2406] = 50'b10_1010110000110000_0111111111010000_0010110000010000;
      patterns[2407] = 50'b11_1010110000110000_0111111111010000_1111111111110000;
      patterns[2408] = 50'b00_1110111000010110_0000111011110110_1111110100001100;
      patterns[2409] = 50'b01_1110111000010110_0000111011110110_1101111100100000;
      patterns[2410] = 50'b10_1110111000010110_0000111011110110_0000111000010110;
      patterns[2411] = 50'b11_1110111000010110_0000111011110110_1110111011110110;
      patterns[2412] = 50'b00_0011111101010100_1000000010101101_1100000000000001;
      patterns[2413] = 50'b01_0011111101010100_1000000010101101_1011111010100111;
      patterns[2414] = 50'b10_0011111101010100_1000000010101101_0000000000000100;
      patterns[2415] = 50'b11_0011111101010100_1000000010101101_1011111111111101;
      patterns[2416] = 50'b00_0011100000110010_1101110111011101_0001011000001111;
      patterns[2417] = 50'b01_0011100000110010_1101110111011101_0101101001010101;
      patterns[2418] = 50'b10_0011100000110010_1101110111011101_0001100000010000;
      patterns[2419] = 50'b11_0011100000110010_1101110111011101_1111110111111111;
      patterns[2420] = 50'b00_0011111100011000_1100101110101110_0000101011000110;
      patterns[2421] = 50'b01_0011111100011000_1100101110101110_0111001101101010;
      patterns[2422] = 50'b10_0011111100011000_1100101110101110_0000101100001000;
      patterns[2423] = 50'b11_0011111100011000_1100101110101110_1111111110111110;
      patterns[2424] = 50'b00_1110001001100000_0101011011001001_0011100100101001;
      patterns[2425] = 50'b01_1110001001100000_0101011011001001_1000101110010111;
      patterns[2426] = 50'b10_1110001001100000_0101011011001001_0100001001000000;
      patterns[2427] = 50'b11_1110001001100000_0101011011001001_1111011011101001;
      patterns[2428] = 50'b00_1001111101010100_1111100100010010_1001100001100110;
      patterns[2429] = 50'b01_1001111101010100_1111100100010010_1010011001000010;
      patterns[2430] = 50'b10_1001111101010100_1111100100010010_1001100100010000;
      patterns[2431] = 50'b11_1001111101010100_1111100100010010_1111111101010110;
      patterns[2432] = 50'b00_0011101110001011_0001010111001101_0101000101011000;
      patterns[2433] = 50'b01_0011101110001011_0001010111001101_0010010110111110;
      patterns[2434] = 50'b10_0011101110001011_0001010111001101_0001000110001001;
      patterns[2435] = 50'b11_0011101110001011_0001010111001101_0011111111001111;
      patterns[2436] = 50'b00_1101000101010010_0000001101001001_1101010010011011;
      patterns[2437] = 50'b01_1101000101010010_0000001101001001_1100111000001001;
      patterns[2438] = 50'b10_1101000101010010_0000001101001001_0000000101000000;
      patterns[2439] = 50'b11_1101000101010010_0000001101001001_1101001101011011;
      patterns[2440] = 50'b00_0100101101000101_0110101000101100_1011010101110001;
      patterns[2441] = 50'b01_0100101101000101_0110101000101100_1110000100011001;
      patterns[2442] = 50'b10_0100101101000101_0110101000101100_0100101000000100;
      patterns[2443] = 50'b11_0100101101000101_0110101000101100_0110101101101101;
      patterns[2444] = 50'b00_1110111110100111_0011010010110010_0010010001011001;
      patterns[2445] = 50'b01_1110111110100111_0011010010110010_1011101011110101;
      patterns[2446] = 50'b10_1110111110100111_0011010010110010_0010010010100010;
      patterns[2447] = 50'b11_1110111110100111_0011010010110010_1111111110110111;
      patterns[2448] = 50'b00_1100011011101010_1101101011101000_1010000111010010;
      patterns[2449] = 50'b01_1100011011101010_1101101011101000_1110110000000010;
      patterns[2450] = 50'b10_1100011011101010_1101101011101000_1100001011101000;
      patterns[2451] = 50'b11_1100011011101010_1101101011101000_1101111011101010;
      patterns[2452] = 50'b00_1010101100010101_1001111101001110_0100101001100011;
      patterns[2453] = 50'b01_1010101100010101_1001111101001110_0000101111000111;
      patterns[2454] = 50'b10_1010101100010101_1001111101001110_1000101100000100;
      patterns[2455] = 50'b11_1010101100010101_1001111101001110_1011111101011111;
      patterns[2456] = 50'b00_0000110100011010_0101000010010011_0101110110101101;
      patterns[2457] = 50'b01_0000110100011010_0101000010010011_1011110010000111;
      patterns[2458] = 50'b10_0000110100011010_0101000010010011_0000000000010010;
      patterns[2459] = 50'b11_0000110100011010_0101000010010011_0101110110011011;
      patterns[2460] = 50'b00_0111001001010001_1001110011001110_0000111100011111;
      patterns[2461] = 50'b01_0111001001010001_1001110011001110_1101010110000011;
      patterns[2462] = 50'b10_0111001001010001_1001110011001110_0001000001000000;
      patterns[2463] = 50'b11_0111001001010001_1001110011001110_1111111011011111;
      patterns[2464] = 50'b00_0010010011110101_1001111101100010_1100010001010111;
      patterns[2465] = 50'b01_0010010011110101_1001111101100010_1000010110010011;
      patterns[2466] = 50'b10_0010010011110101_1001111101100010_0000010001100000;
      patterns[2467] = 50'b11_0010010011110101_1001111101100010_1011111111110111;
      patterns[2468] = 50'b00_1110111111001000_0111100010100110_0110100001101110;
      patterns[2469] = 50'b01_1110111111001000_0111100010100110_0111011100100010;
      patterns[2470] = 50'b10_1110111111001000_0111100010100110_0110100010000000;
      patterns[2471] = 50'b11_1110111111001000_0111100010100110_1111111111101110;
      patterns[2472] = 50'b00_0011001111011011_1100001111011101_1111011110111000;
      patterns[2473] = 50'b01_0011001111011011_1100001111011101_0110111111111110;
      patterns[2474] = 50'b10_0011001111011011_1100001111011101_0000001111011001;
      patterns[2475] = 50'b11_0011001111011011_1100001111011101_1111001111011111;
      patterns[2476] = 50'b00_1000000110111100_0011000100010011_1011001011001111;
      patterns[2477] = 50'b01_1000000110111100_0011000100010011_0101000010101001;
      patterns[2478] = 50'b10_1000000110111100_0011000100010011_0000000100010000;
      patterns[2479] = 50'b11_1000000110111100_0011000100010011_1011000110111111;
      patterns[2480] = 50'b00_1011100110100110_0110001110100001_0001110101000111;
      patterns[2481] = 50'b01_1011100110100110_0110001110100001_0101011000000101;
      patterns[2482] = 50'b10_1011100110100110_0110001110100001_0010000110100000;
      patterns[2483] = 50'b11_1011100110100110_0110001110100001_1111101110100111;
      patterns[2484] = 50'b00_1100001001001001_0010111100110011_1111000101111100;
      patterns[2485] = 50'b01_1100001001001001_0010111100110011_1001001100010110;
      patterns[2486] = 50'b10_1100001001001001_0010111100110011_0000001000000001;
      patterns[2487] = 50'b11_1100001001001001_0010111100110011_1110111101111011;
      patterns[2488] = 50'b00_0010100010100011_0000101100010000_0011001110110011;
      patterns[2489] = 50'b01_0010100010100011_0000101100010000_0001110110010011;
      patterns[2490] = 50'b10_0010100010100011_0000101100010000_0000100000000000;
      patterns[2491] = 50'b11_0010100010100011_0000101100010000_0010101110110011;
      patterns[2492] = 50'b00_1000111001000111_1111000110101001_0111111111110000;
      patterns[2493] = 50'b01_1000111001000111_1111000110101001_1001110010011110;
      patterns[2494] = 50'b10_1000111001000111_1111000110101001_1000000000000001;
      patterns[2495] = 50'b11_1000111001000111_1111000110101001_1111111111101111;
      patterns[2496] = 50'b00_0001101110101111_0010111111110000_0100101110011111;
      patterns[2497] = 50'b01_0001101110101111_0010111111110000_1110101110111111;
      patterns[2498] = 50'b10_0001101110101111_0010111111110000_0000101110100000;
      patterns[2499] = 50'b11_0001101110101111_0010111111110000_0011111111111111;
      patterns[2500] = 50'b00_0011101011111110_1110100001101111_0010001101101101;
      patterns[2501] = 50'b01_0011101011111110_1110100001101111_0101001010001111;
      patterns[2502] = 50'b10_0011101011111110_1110100001101111_0010100001101110;
      patterns[2503] = 50'b11_0011101011111110_1110100001101111_1111101011111111;
      patterns[2504] = 50'b00_1000001001000111_0011100001000101_1011101010001100;
      patterns[2505] = 50'b01_1000001001000111_0011100001000101_0100101000000010;
      patterns[2506] = 50'b10_1000001001000111_0011100001000101_0000000001000101;
      patterns[2507] = 50'b11_1000001001000111_0011100001000101_1011101001000111;
      patterns[2508] = 50'b00_1101010000100110_0010101110110110_1111111111011100;
      patterns[2509] = 50'b01_1101010000100110_0010101110110110_1010100001110000;
      patterns[2510] = 50'b10_1101010000100110_0010101110110110_0000000000100110;
      patterns[2511] = 50'b11_1101010000100110_0010101110110110_1111111110110110;
      patterns[2512] = 50'b00_1001011101111001_1010001111101011_0011101101100100;
      patterns[2513] = 50'b01_1001011101111001_1010001111101011_1111001110001110;
      patterns[2514] = 50'b10_1001011101111001_1010001111101011_1000001101101001;
      patterns[2515] = 50'b11_1001011101111001_1010001111101011_1011011111111011;
      patterns[2516] = 50'b00_0100110010111101_0100101100010100_1001011111010001;
      patterns[2517] = 50'b01_0100110010111101_0100101100010100_0000000110101001;
      patterns[2518] = 50'b10_0100110010111101_0100101100010100_0100100000010100;
      patterns[2519] = 50'b11_0100110010111101_0100101100010100_0100111110111101;
      patterns[2520] = 50'b00_0101110111110100_1111111011001010_0101110010111110;
      patterns[2521] = 50'b01_0101110111110100_1111111011001010_0101111100101010;
      patterns[2522] = 50'b10_0101110111110100_1111111011001010_0101110011000000;
      patterns[2523] = 50'b11_0101110111110100_1111111011001010_1111111111111110;
      patterns[2524] = 50'b00_1000011010001111_0010110101010100_1011001111100011;
      patterns[2525] = 50'b01_1000011010001111_0010110101010100_0101100100111011;
      patterns[2526] = 50'b10_1000011010001111_0010110101010100_0000010000000100;
      patterns[2527] = 50'b11_1000011010001111_0010110101010100_1010111111011111;
      patterns[2528] = 50'b00_1010100010110001_0111000010010111_0001100101001000;
      patterns[2529] = 50'b01_1010100010110001_0111000010010111_0011100000011010;
      patterns[2530] = 50'b10_1010100010110001_0111000010010111_0010000010010001;
      patterns[2531] = 50'b11_1010100010110001_0111000010010111_1111100010110111;
      patterns[2532] = 50'b00_1111010110001101_1101110010100100_1101001000110001;
      patterns[2533] = 50'b01_1111010110001101_1101110010100100_0001100011101001;
      patterns[2534] = 50'b10_1111010110001101_1101110010100100_1101010010000100;
      patterns[2535] = 50'b11_1111010110001101_1101110010100100_1111110110101101;
      patterns[2536] = 50'b00_0110110011101101_1001011001111110_0000001101101011;
      patterns[2537] = 50'b01_0110110011101101_1001011001111110_1101011001101111;
      patterns[2538] = 50'b10_0110110011101101_1001011001111110_0000010001101100;
      patterns[2539] = 50'b11_0110110011101101_1001011001111110_1111111011111111;
      patterns[2540] = 50'b00_0110110101000111_0010010111111110_1001001101000101;
      patterns[2541] = 50'b01_0110110101000111_0010010111111110_0100011101001001;
      patterns[2542] = 50'b10_0110110101000111_0010010111111110_0010010101000110;
      patterns[2543] = 50'b11_0110110101000111_0010010111111110_0110110111111111;
      patterns[2544] = 50'b00_0011011101101111_1101001000110110_0000100110100101;
      patterns[2545] = 50'b01_0011011101101111_1101001000110110_0110010100111001;
      patterns[2546] = 50'b10_0011011101101111_1101001000110110_0001001000100110;
      patterns[2547] = 50'b11_0011011101101111_1101001000110110_1111011101111111;
      patterns[2548] = 50'b00_0101100000110010_0010010111110111_0111111000101001;
      patterns[2549] = 50'b01_0101100000110010_0010010111110111_0011001000111011;
      patterns[2550] = 50'b10_0101100000110010_0010010111110111_0000000000110010;
      patterns[2551] = 50'b11_0101100000110010_0010010111110111_0111110111110111;
      patterns[2552] = 50'b00_0010010001010111_0110000101010010_1000010110101001;
      patterns[2553] = 50'b01_0010010001010111_0110000101010010_1100001100000101;
      patterns[2554] = 50'b10_0010010001010111_0110000101010010_0010000001010010;
      patterns[2555] = 50'b11_0010010001010111_0110000101010010_0110010101010111;
      patterns[2556] = 50'b00_0011000101111010_0011100001101110_0110100111101000;
      patterns[2557] = 50'b01_0011000101111010_0011100001101110_1111100100001100;
      patterns[2558] = 50'b10_0011000101111010_0011100001101110_0011000001101010;
      patterns[2559] = 50'b11_0011000101111010_0011100001101110_0011100101111110;
      patterns[2560] = 50'b00_1010010111101010_0101111011001000_0000010010110010;
      patterns[2561] = 50'b01_1010010111101010_0101111011001000_0100011100100010;
      patterns[2562] = 50'b10_1010010111101010_0101111011001000_0000010011001000;
      patterns[2563] = 50'b11_1010010111101010_0101111011001000_1111111111101010;
      patterns[2564] = 50'b00_1001101110010110_0100001110101011_1101111101000001;
      patterns[2565] = 50'b01_1001101110010110_0100001110101011_0101011111101011;
      patterns[2566] = 50'b10_1001101110010110_0100001110101011_0000001110000010;
      patterns[2567] = 50'b11_1001101110010110_0100001110101011_1101101110111111;
      patterns[2568] = 50'b00_1011110000011011_0100100000001111_0000010000101010;
      patterns[2569] = 50'b01_1011110000011011_0100100000001111_0111010000001100;
      patterns[2570] = 50'b10_1011110000011011_0100100000001111_0000100000001011;
      patterns[2571] = 50'b11_1011110000011011_0100100000001111_1111110000011111;
      patterns[2572] = 50'b00_1101011011101000_0000001011110010_1101100111011010;
      patterns[2573] = 50'b01_1101011011101000_0000001011110010_1101001111110110;
      patterns[2574] = 50'b10_1101011011101000_0000001011110010_0000001011100000;
      patterns[2575] = 50'b11_1101011011101000_0000001011110010_1101011011111010;
      patterns[2576] = 50'b00_1111101111000111_1011111001000111_1011101000001110;
      patterns[2577] = 50'b01_1111101111000111_1011111001000111_0011110110000000;
      patterns[2578] = 50'b10_1111101111000111_1011111001000111_1011101001000111;
      patterns[2579] = 50'b11_1111101111000111_1011111001000111_1111111111000111;
      patterns[2580] = 50'b00_1010110011111111_1100011110011011_0111010010011010;
      patterns[2581] = 50'b01_1010110011111111_1100011110011011_1110010101100100;
      patterns[2582] = 50'b10_1010110011111111_1100011110011011_1000010010011011;
      patterns[2583] = 50'b11_1010110011111111_1100011110011011_1110111111111111;
      patterns[2584] = 50'b00_1110100111011111_0000001101000110_1110110100100101;
      patterns[2585] = 50'b01_1110100111011111_0000001101000110_1110011010011001;
      patterns[2586] = 50'b10_1110100111011111_0000001101000110_0000000101000110;
      patterns[2587] = 50'b11_1110100111011111_0000001101000110_1110101111011111;
      patterns[2588] = 50'b00_0001111001101011_0010001100110010_0100000110011101;
      patterns[2589] = 50'b01_0001111001101011_0010001100110010_1111101100111001;
      patterns[2590] = 50'b10_0001111001101011_0010001100110010_0000001000100010;
      patterns[2591] = 50'b11_0001111001101011_0010001100110010_0011111101111011;
      patterns[2592] = 50'b00_1011101111111001_0010000110001111_1101110110001000;
      patterns[2593] = 50'b01_1011101111111001_0010000110001111_1001101001101010;
      patterns[2594] = 50'b10_1011101111111001_0010000110001111_0010000110001001;
      patterns[2595] = 50'b11_1011101111111001_0010000110001111_1011101111111111;
      patterns[2596] = 50'b00_0100001000011101_0001000000110111_0101001001010100;
      patterns[2597] = 50'b01_0100001000011101_0001000000110111_0011000111100110;
      patterns[2598] = 50'b10_0100001000011101_0001000000110111_0000000000010101;
      patterns[2599] = 50'b11_0100001000011101_0001000000110111_0101001000111111;
      patterns[2600] = 50'b00_1000010100001001_1100010101110101_0100101001111110;
      patterns[2601] = 50'b01_1000010100001001_1100010101110101_1011111110010100;
      patterns[2602] = 50'b10_1000010100001001_1100010101110101_1000010100000001;
      patterns[2603] = 50'b11_1000010100001001_1100010101110101_1100010101111101;
      patterns[2604] = 50'b00_1100111011001110_0111101001101011_0100100100111001;
      patterns[2605] = 50'b01_1100111011001110_0111101001101011_0101010001100011;
      patterns[2606] = 50'b10_1100111011001110_0111101001101011_0100101001001010;
      patterns[2607] = 50'b11_1100111011001110_0111101001101011_1111111011101111;
      patterns[2608] = 50'b00_0011001000110000_1000110100000010_1011111100110010;
      patterns[2609] = 50'b01_0011001000110000_1000110100000010_1010010100101110;
      patterns[2610] = 50'b10_0011001000110000_1000110100000010_0000000000000000;
      patterns[2611] = 50'b11_0011001000110000_1000110100000010_1011111100110010;
      patterns[2612] = 50'b00_1011011111101011_0111101011100000_0011001011001011;
      patterns[2613] = 50'b01_1011011111101011_0111101011100000_0011110100001011;
      patterns[2614] = 50'b10_1011011111101011_0111101011100000_0011001011100000;
      patterns[2615] = 50'b11_1011011111101011_0111101011100000_1111111111101011;
      patterns[2616] = 50'b00_1000000011100011_1111101101100010_0111110001000101;
      patterns[2617] = 50'b01_1000000011100011_1111101101100010_1000010110000001;
      patterns[2618] = 50'b10_1000000011100011_1111101101100010_1000000001100010;
      patterns[2619] = 50'b11_1000000011100011_1111101101100010_1111101111100011;
      patterns[2620] = 50'b00_0010000011110100_0011011100100001_0101100000010101;
      patterns[2621] = 50'b01_0010000011110100_0011011100100001_1110100111010011;
      patterns[2622] = 50'b10_0010000011110100_0011011100100001_0010000000100000;
      patterns[2623] = 50'b11_0010000011110100_0011011100100001_0011011111110101;
      patterns[2624] = 50'b00_0100010011100110_0100101111011011_1001000011000001;
      patterns[2625] = 50'b01_0100010011100110_0100101111011011_1111100100001011;
      patterns[2626] = 50'b10_0100010011100110_0100101111011011_0100000011000010;
      patterns[2627] = 50'b11_0100010011100110_0100101111011011_0100111111111111;
      patterns[2628] = 50'b00_1010101101100001_0001011000110001_1100000110010010;
      patterns[2629] = 50'b01_1010101101100001_0001011000110001_1001010100110000;
      patterns[2630] = 50'b10_1010101101100001_0001011000110001_0000001000100001;
      patterns[2631] = 50'b11_1010101101100001_0001011000110001_1011111101110001;
      patterns[2632] = 50'b00_1110100111001100_0001011110101001_0000000101110101;
      patterns[2633] = 50'b01_1110100111001100_0001011110101001_1101001000100011;
      patterns[2634] = 50'b10_1110100111001100_0001011110101001_0000000110001000;
      patterns[2635] = 50'b11_1110100111001100_0001011110101001_1111111111101101;
      patterns[2636] = 50'b00_1100110001011100_1110100100111101_1011010110011001;
      patterns[2637] = 50'b01_1100110001011100_1110100100111101_1110001100011111;
      patterns[2638] = 50'b10_1100110001011100_1110100100111101_1100100000011100;
      patterns[2639] = 50'b11_1100110001011100_1110100100111101_1110110101111101;
      patterns[2640] = 50'b00_0001100011111100_0010000100110101_0011101000110001;
      patterns[2641] = 50'b01_0001100011111100_0010000100110101_1111011111000111;
      patterns[2642] = 50'b10_0001100011111100_0010000100110101_0000000000110100;
      patterns[2643] = 50'b11_0001100011111100_0010000100110101_0011100111111101;
      patterns[2644] = 50'b00_0110100100000010_1011100100110110_0010001000111000;
      patterns[2645] = 50'b01_0110100100000010_1011100100110110_1010111111001100;
      patterns[2646] = 50'b10_0110100100000010_1011100100110110_0010100100000010;
      patterns[2647] = 50'b11_0110100100000010_1011100100110110_1111100100110110;
      patterns[2648] = 50'b00_1101001001111010_1001111010000001_0111000011111011;
      patterns[2649] = 50'b01_1101001001111010_1001111010000001_0011001111111001;
      patterns[2650] = 50'b10_1101001001111010_1001111010000001_1001001000000000;
      patterns[2651] = 50'b11_1101001001111010_1001111010000001_1101111011111011;
      patterns[2652] = 50'b00_0111000011101110_0010010110101011_1001011010011001;
      patterns[2653] = 50'b01_0111000011101110_0010010110101011_0100101101000011;
      patterns[2654] = 50'b10_0111000011101110_0010010110101011_0010000010101010;
      patterns[2655] = 50'b11_0111000011101110_0010010110101011_0111010111101111;
      patterns[2656] = 50'b00_0001001111100001_0000101111001011_0001111110101100;
      patterns[2657] = 50'b01_0001001111100001_0000101111001011_0000100000010110;
      patterns[2658] = 50'b10_0001001111100001_0000101111001011_0000001111000001;
      patterns[2659] = 50'b11_0001001111100001_0000101111001011_0001101111101011;
      patterns[2660] = 50'b00_1001000000110100_1010010010100110_0011010011011010;
      patterns[2661] = 50'b01_1001000000110100_1010010010100110_1110101110001110;
      patterns[2662] = 50'b10_1001000000110100_1010010010100110_1000000000100100;
      patterns[2663] = 50'b11_1001000000110100_1010010010100110_1011010010110110;
      patterns[2664] = 50'b00_0101111001010111_1110011010101111_0100010100000110;
      patterns[2665] = 50'b01_0101111001010111_1110011010101111_0111011110101000;
      patterns[2666] = 50'b10_0101111001010111_1110011010101111_0100011000000111;
      patterns[2667] = 50'b11_0101111001010111_1110011010101111_1111111011111111;
      patterns[2668] = 50'b00_0101101100100110_0111111001011111_1101100110000101;
      patterns[2669] = 50'b01_0101101100100110_0111111001011111_1101110011000111;
      patterns[2670] = 50'b10_0101101100100110_0111111001011111_0101101000000110;
      patterns[2671] = 50'b11_0101101100100110_0111111001011111_0111111101111111;
      patterns[2672] = 50'b00_0000100101100010_1011000101100010_1011101011000100;
      patterns[2673] = 50'b01_0000100101100010_1011000101100010_0101100000000000;
      patterns[2674] = 50'b10_0000100101100010_1011000101100010_0000000101100010;
      patterns[2675] = 50'b11_0000100101100010_1011000101100010_1011100101100010;
      patterns[2676] = 50'b00_1000011101110101_0001001100000000_1001101001110101;
      patterns[2677] = 50'b01_1000011101110101_0001001100000000_0111010001110101;
      patterns[2678] = 50'b10_1000011101110101_0001001100000000_0000001100000000;
      patterns[2679] = 50'b11_1000011101110101_0001001100000000_1001011101110101;
      patterns[2680] = 50'b00_0101010111101111_0100010010110010_1001101010100001;
      patterns[2681] = 50'b01_0101010111101111_0100010010110010_0001000100111101;
      patterns[2682] = 50'b10_0101010111101111_0100010010110010_0100010010100010;
      patterns[2683] = 50'b11_0101010111101111_0100010010110010_0101010111111111;
      patterns[2684] = 50'b00_1101111110010000_1101001111011001_1011001101101001;
      patterns[2685] = 50'b01_1101111110010000_1101001111011001_0000101110110111;
      patterns[2686] = 50'b10_1101111110010000_1101001111011001_1101001110010000;
      patterns[2687] = 50'b11_1101111110010000_1101001111011001_1101111111011001;
      patterns[2688] = 50'b00_1010000111110110_1100011011110101_0110100011101011;
      patterns[2689] = 50'b01_1010000111110110_1100011011110101_1101101100000001;
      patterns[2690] = 50'b10_1010000111110110_1100011011110101_1000000011110100;
      patterns[2691] = 50'b11_1010000111110110_1100011011110101_1110011111110111;
      patterns[2692] = 50'b00_1001111001011100_0101110010101101_1111101100001001;
      patterns[2693] = 50'b01_1001111001011100_0101110010101101_0100000110101111;
      patterns[2694] = 50'b10_1001111001011100_0101110010101101_0001110000001100;
      patterns[2695] = 50'b11_1001111001011100_0101110010101101_1101111011111101;
      patterns[2696] = 50'b00_1111001001110001_1001010100011110_1000011110001111;
      patterns[2697] = 50'b01_1111001001110001_1001010100011110_0101110101010011;
      patterns[2698] = 50'b10_1111001001110001_1001010100011110_1001000000010000;
      patterns[2699] = 50'b11_1111001001110001_1001010100011110_1111011101111111;
      patterns[2700] = 50'b00_1100101010010010_0100010100010101_0000111110100111;
      patterns[2701] = 50'b01_1100101010010010_0100010100010101_1000010101111101;
      patterns[2702] = 50'b10_1100101010010010_0100010100010101_0100000000010000;
      patterns[2703] = 50'b11_1100101010010010_0100010100010101_1100111110010111;
      patterns[2704] = 50'b00_0100011010110010_0000101010000111_0101000100111001;
      patterns[2705] = 50'b01_0100011010110010_0000101010000111_0011110000101011;
      patterns[2706] = 50'b10_0100011010110010_0000101010000111_0000001010000010;
      patterns[2707] = 50'b11_0100011010110010_0000101010000111_0100111010110111;
      patterns[2708] = 50'b00_1111101001110011_1001010100000101_1000111101111000;
      patterns[2709] = 50'b01_1111101001110011_1001010100000101_0110010101101110;
      patterns[2710] = 50'b10_1111101001110011_1001010100000101_1001000000000001;
      patterns[2711] = 50'b11_1111101001110011_1001010100000101_1111111101110111;
      patterns[2712] = 50'b00_1100110101000010_0101101100110110_0010100001111000;
      patterns[2713] = 50'b01_1100110101000010_0101101100110110_0111001000001100;
      patterns[2714] = 50'b10_1100110101000010_0101101100110110_0100100100000010;
      patterns[2715] = 50'b11_1100110101000010_0101101100110110_1101111101110110;
      patterns[2716] = 50'b00_1010000110010001_0100001011110110_1110010010000111;
      patterns[2717] = 50'b01_1010000110010001_0100001011110110_0101111010011011;
      patterns[2718] = 50'b10_1010000110010001_0100001011110110_0000000010010000;
      patterns[2719] = 50'b11_1010000110010001_0100001011110110_1110001111110111;
      patterns[2720] = 50'b00_0001111111000111_1010001110110011_1100001101111010;
      patterns[2721] = 50'b01_0001111111000111_1010001110110011_0111110000010100;
      patterns[2722] = 50'b10_0001111111000111_1010001110110011_0000001110000011;
      patterns[2723] = 50'b11_0001111111000111_1010001110110011_1011111111110111;
      patterns[2724] = 50'b00_1010101111100100_1100010101010101_0111000100111001;
      patterns[2725] = 50'b01_1010101111100100_1100010101010101_1110011010001111;
      patterns[2726] = 50'b10_1010101111100100_1100010101010101_1000000101000100;
      patterns[2727] = 50'b11_1010101111100100_1100010101010101_1110111111110101;
      patterns[2728] = 50'b00_0010000010101110_1110100010101001_0000100101010111;
      patterns[2729] = 50'b01_0010000010101110_1110100010101001_0011100000000101;
      patterns[2730] = 50'b10_0010000010101110_1110100010101001_0010000010101000;
      patterns[2731] = 50'b11_0010000010101110_1110100010101001_1110100010101111;
      patterns[2732] = 50'b00_1011001001101010_1000110000011110_0011111010001000;
      patterns[2733] = 50'b01_1011001001101010_1000110000011110_0010011001001100;
      patterns[2734] = 50'b10_1011001001101010_1000110000011110_1000000000001010;
      patterns[2735] = 50'b11_1011001001101010_1000110000011110_1011111001111110;
      patterns[2736] = 50'b00_1111001010010100_1111111111101010_1111001001111110;
      patterns[2737] = 50'b01_1111001010010100_1111111111101010_1111001010101010;
      patterns[2738] = 50'b10_1111001010010100_1111111111101010_1111001010000000;
      patterns[2739] = 50'b11_1111001010010100_1111111111101010_1111111111111110;
      patterns[2740] = 50'b00_1000011011111101_0010101011010100_1011000111010001;
      patterns[2741] = 50'b01_1000011011111101_0010101011010100_0101110000101001;
      patterns[2742] = 50'b10_1000011011111101_0010101011010100_0000001011010100;
      patterns[2743] = 50'b11_1000011011111101_0010101011010100_1010111011111101;
      patterns[2744] = 50'b00_1100011010011110_0100001110010100_0000101000110010;
      patterns[2745] = 50'b01_1100011010011110_0100001110010100_1000001100001010;
      patterns[2746] = 50'b10_1100011010011110_0100001110010100_0100001010010100;
      patterns[2747] = 50'b11_1100011010011110_0100001110010100_1100011110011110;
      patterns[2748] = 50'b00_0010111000111001_0001011000111101_0100010001110110;
      patterns[2749] = 50'b01_0010111000111001_0001011000111101_0001011111111100;
      patterns[2750] = 50'b10_0010111000111001_0001011000111101_0000011000111001;
      patterns[2751] = 50'b11_0010111000111001_0001011000111101_0011111000111101;
      patterns[2752] = 50'b00_1110110001001101_0111111101101010_0110101110110111;
      patterns[2753] = 50'b01_1110110001001101_0111111101101010_0110110011100011;
      patterns[2754] = 50'b10_1110110001001101_0111111101101010_0110110001001000;
      patterns[2755] = 50'b11_1110110001001101_0111111101101010_1111111101101111;
      patterns[2756] = 50'b00_1001111101111111_0001110010001010_1011110000001001;
      patterns[2757] = 50'b01_1001111101111111_0001110010001010_1000001011110101;
      patterns[2758] = 50'b10_1001111101111111_0001110010001010_0001110000001010;
      patterns[2759] = 50'b11_1001111101111111_0001110010001010_1001111111111111;
      patterns[2760] = 50'b00_1010001001101110_1011111110101011_0110001000011001;
      patterns[2761] = 50'b01_1010001001101110_1011111110101011_1110001011000011;
      patterns[2762] = 50'b10_1010001001101110_1011111110101011_1010001000101010;
      patterns[2763] = 50'b11_1010001001101110_1011111110101011_1011111111101111;
      patterns[2764] = 50'b00_1100110001111100_0010100111011000_1111011001010100;
      patterns[2765] = 50'b01_1100110001111100_0010100111011000_1010001010100100;
      patterns[2766] = 50'b10_1100110001111100_0010100111011000_0000100001011000;
      patterns[2767] = 50'b11_1100110001111100_0010100111011000_1110110111111100;
      patterns[2768] = 50'b00_1010011000111100_1000011111100100_0010111000100000;
      patterns[2769] = 50'b01_1010011000111100_1000011111100100_0001111001011000;
      patterns[2770] = 50'b10_1010011000111100_1000011111100100_1000011000100100;
      patterns[2771] = 50'b11_1010011000111100_1000011111100100_1010011111111100;
      patterns[2772] = 50'b00_1000001011001010_0111111000110001_0000000011111011;
      patterns[2773] = 50'b01_1000001011001010_0111111000110001_0000010010011001;
      patterns[2774] = 50'b10_1000001011001010_0111111000110001_0000001000000000;
      patterns[2775] = 50'b11_1000001011001010_0111111000110001_1111111011111011;
      patterns[2776] = 50'b00_0110001011010011_0111111110011101_1110001001110000;
      patterns[2777] = 50'b01_0110001011010011_0111111110011101_1110001100110110;
      patterns[2778] = 50'b10_0110001011010011_0111111110011101_0110001010010001;
      patterns[2779] = 50'b11_0110001011010011_0111111110011101_0111111111011111;
      patterns[2780] = 50'b00_1011001110000010_0011010101111101_1110100011111111;
      patterns[2781] = 50'b01_1011001110000010_0011010101111101_0111111000000101;
      patterns[2782] = 50'b10_1011001110000010_0011010101111101_0011000100000000;
      patterns[2783] = 50'b11_1011001110000010_0011010101111101_1011011111111111;
      patterns[2784] = 50'b00_1111000010001010_1101000111011000_1100001001100010;
      patterns[2785] = 50'b01_1111000010001010_1101000111011000_0001111010110010;
      patterns[2786] = 50'b10_1111000010001010_1101000111011000_1101000010001000;
      patterns[2787] = 50'b11_1111000010001010_1101000111011000_1111000111011010;
      patterns[2788] = 50'b00_1000110111011010_1110010100000011_0111001011011101;
      patterns[2789] = 50'b01_1000110111011010_1110010100000011_1010100011010111;
      patterns[2790] = 50'b10_1000110111011010_1110010100000011_1000010100000010;
      patterns[2791] = 50'b11_1000110111011010_1110010100000011_1110110111011011;
      patterns[2792] = 50'b00_1100100011010010_0101001110101110_0001110010000000;
      patterns[2793] = 50'b01_1100100011010010_0101001110101110_0111010100100100;
      patterns[2794] = 50'b10_1100100011010010_0101001110101110_0100000010000010;
      patterns[2795] = 50'b11_1100100011010010_0101001110101110_1101101111111110;
      patterns[2796] = 50'b00_1010001100110011_0001110101110000_1100000010100011;
      patterns[2797] = 50'b01_1010001100110011_0001110101110000_1000010111000011;
      patterns[2798] = 50'b10_1010001100110011_0001110101110000_0000000100110000;
      patterns[2799] = 50'b11_1010001100110011_0001110101110000_1011111101110011;
      patterns[2800] = 50'b00_0011000010101001_0000010110100111_0011011001010000;
      patterns[2801] = 50'b01_0011000010101001_0000010110100111_0010101100000010;
      patterns[2802] = 50'b10_0011000010101001_0000010110100111_0000000010100001;
      patterns[2803] = 50'b11_0011000010101001_0000010110100111_0011010110101111;
      patterns[2804] = 50'b00_1111110000011000_1101001110000001_1100111110011001;
      patterns[2805] = 50'b01_1111110000011000_1101001110000001_0010100010010111;
      patterns[2806] = 50'b10_1111110000011000_1101001110000001_1101000000000000;
      patterns[2807] = 50'b11_1111110000011000_1101001110000001_1111111110011001;
      patterns[2808] = 50'b00_1110000011010001_1010101001111010_1000101101001011;
      patterns[2809] = 50'b01_1110000011010001_1010101001111010_0011011001010111;
      patterns[2810] = 50'b10_1110000011010001_1010101001111010_1010000001010000;
      patterns[2811] = 50'b11_1110000011010001_1010101001111010_1110101011111011;
      patterns[2812] = 50'b00_1001111100101100_0000110011001001_1010101111110101;
      patterns[2813] = 50'b01_1001111100101100_0000110011001001_1001001001100011;
      patterns[2814] = 50'b10_1001111100101100_0000110011001001_0000110000001000;
      patterns[2815] = 50'b11_1001111100101100_0000110011001001_1001111111101101;
      patterns[2816] = 50'b00_0110000001001000_1111110101010111_0101110110011111;
      patterns[2817] = 50'b01_0110000001001000_1111110101010111_0110001011110001;
      patterns[2818] = 50'b10_0110000001001000_1111110101010111_0110000001000000;
      patterns[2819] = 50'b11_0110000001001000_1111110101010111_1111110101011111;
      patterns[2820] = 50'b00_1000101111111100_1011000100101100_0011110100101000;
      patterns[2821] = 50'b01_1000101111111100_1011000100101100_1101101011010000;
      patterns[2822] = 50'b10_1000101111111100_1011000100101100_1000000100101100;
      patterns[2823] = 50'b11_1000101111111100_1011000100101100_1011101111111100;
      patterns[2824] = 50'b00_1101101010111000_1000100011111001_0110001110110001;
      patterns[2825] = 50'b01_1101101010111000_1000100011111001_0101000110111111;
      patterns[2826] = 50'b10_1101101010111000_1000100011111001_1000100010111000;
      patterns[2827] = 50'b11_1101101010111000_1000100011111001_1101101011111001;
      patterns[2828] = 50'b00_1001010100101101_0000110100001000_1010001000110101;
      patterns[2829] = 50'b01_1001010100101101_0000110100001000_1000100000100101;
      patterns[2830] = 50'b10_1001010100101101_0000110100001000_0000010100001000;
      patterns[2831] = 50'b11_1001010100101101_0000110100001000_1001110100101101;
      patterns[2832] = 50'b00_1111100111011111_0100000000001011_0011100111101010;
      patterns[2833] = 50'b01_1111100111011111_0100000000001011_1011100111010100;
      patterns[2834] = 50'b10_1111100111011111_0100000000001011_0100000000001011;
      patterns[2835] = 50'b11_1111100111011111_0100000000001011_1111100111011111;
      patterns[2836] = 50'b00_1101011010001010_0110001100110000_0011100110111010;
      patterns[2837] = 50'b01_1101011010001010_0110001100110000_0111001101011010;
      patterns[2838] = 50'b10_1101011010001010_0110001100110000_0100001000000000;
      patterns[2839] = 50'b11_1101011010001010_0110001100110000_1111011110111010;
      patterns[2840] = 50'b00_0110111000100011_1011111010110000_0010110011010011;
      patterns[2841] = 50'b01_0110111000100011_1011111010110000_1010111101110011;
      patterns[2842] = 50'b10_0110111000100011_1011111010110000_0010111000100000;
      patterns[2843] = 50'b11_0110111000100011_1011111010110000_1111111010110011;
      patterns[2844] = 50'b00_1011110011011100_1110100100011101_1010010111111001;
      patterns[2845] = 50'b01_1011110011011100_1110100100011101_1101001110111111;
      patterns[2846] = 50'b10_1011110011011100_1110100100011101_1010100000011100;
      patterns[2847] = 50'b11_1011110011011100_1110100100011101_1111110111011101;
      patterns[2848] = 50'b00_0101111111010000_1000110000101111_1110101111111111;
      patterns[2849] = 50'b01_0101111111010000_1000110000101111_1101001110100001;
      patterns[2850] = 50'b10_0101111111010000_1000110000101111_0000110000000000;
      patterns[2851] = 50'b11_0101111111010000_1000110000101111_1101111111111111;
      patterns[2852] = 50'b00_1011011010011100_1010101100001011_0110000110100111;
      patterns[2853] = 50'b01_1011011010011100_1010101100001011_0000101110010001;
      patterns[2854] = 50'b10_1011011010011100_1010101100001011_1010001000001000;
      patterns[2855] = 50'b11_1011011010011100_1010101100001011_1011111110011111;
      patterns[2856] = 50'b00_1111011110110011_1100101100010111_1100001011001010;
      patterns[2857] = 50'b01_1111011110110011_1100101100010111_0010110010011100;
      patterns[2858] = 50'b10_1111011110110011_1100101100010111_1100001100010011;
      patterns[2859] = 50'b11_1111011110110011_1100101100010111_1111111110110111;
      patterns[2860] = 50'b00_1010110111011011_0010000011100010_1100111010111101;
      patterns[2861] = 50'b01_1010110111011011_0010000011100010_1000110011111001;
      patterns[2862] = 50'b10_1010110111011011_0010000011100010_0010000011000010;
      patterns[2863] = 50'b11_1010110111011011_0010000011100010_1010110111111011;
      patterns[2864] = 50'b00_1000101100011011_1000010101011010_0001000001110101;
      patterns[2865] = 50'b01_1000101100011011_1000010101011010_0000010111000001;
      patterns[2866] = 50'b10_1000101100011011_1000010101011010_1000000100011010;
      patterns[2867] = 50'b11_1000101100011011_1000010101011010_1000111101011011;
      patterns[2868] = 50'b00_0101110100000011_1011000000011100_0000110100011111;
      patterns[2869] = 50'b01_0101110100000011_1011000000011100_1010110011100111;
      patterns[2870] = 50'b10_0101110100000011_1011000000011100_0001000000000000;
      patterns[2871] = 50'b11_0101110100000011_1011000000011100_1111110100011111;
      patterns[2872] = 50'b00_1011110001100111_0010100100110011_1110010110011010;
      patterns[2873] = 50'b01_1011110001100111_0010100100110011_1001001100110100;
      patterns[2874] = 50'b10_1011110001100111_0010100100110011_0010100000100011;
      patterns[2875] = 50'b11_1011110001100111_0010100100110011_1011110101110111;
      patterns[2876] = 50'b00_0110100100110101_1111001000001100_0101101101000001;
      patterns[2877] = 50'b01_0110100100110101_1111001000001100_0111011100101001;
      patterns[2878] = 50'b10_0110100100110101_1111001000001100_0110000000000100;
      patterns[2879] = 50'b11_0110100100110101_1111001000001100_1111101100111101;
      patterns[2880] = 50'b00_0000111010100110_1101101011011101_1110100110000011;
      patterns[2881] = 50'b01_0000111010100110_1101101011011101_0011001111001001;
      patterns[2882] = 50'b10_0000111010100110_1101101011011101_0000101010000100;
      patterns[2883] = 50'b11_0000111010100110_1101101011011101_1101111011111111;
      patterns[2884] = 50'b00_1110111001111101_0101100100110010_0100011110101111;
      patterns[2885] = 50'b01_1110111001111101_0101100100110010_1001010101001011;
      patterns[2886] = 50'b10_1110111001111101_0101100100110010_0100100000110000;
      patterns[2887] = 50'b11_1110111001111101_0101100100110010_1111111101111111;
      patterns[2888] = 50'b00_0000000000001100_1111011001100011_1111011001101111;
      patterns[2889] = 50'b01_0000000000001100_1111011001100011_0000100110101001;
      patterns[2890] = 50'b10_0000000000001100_1111011001100011_0000000000000000;
      patterns[2891] = 50'b11_0000000000001100_1111011001100011_1111011001101111;
      patterns[2892] = 50'b00_1101001100011000_1011101110001011_1000111010100011;
      patterns[2893] = 50'b01_1101001100011000_1011101110001011_0001011110001101;
      patterns[2894] = 50'b10_1101001100011000_1011101110001011_1001001100001000;
      patterns[2895] = 50'b11_1101001100011000_1011101110001011_1111101110011011;
      patterns[2896] = 50'b00_1011110000010111_0111110000010011_0011100000101010;
      patterns[2897] = 50'b01_1011110000010111_0111110000010011_0100000000000100;
      patterns[2898] = 50'b10_1011110000010111_0111110000010011_0011110000010011;
      patterns[2899] = 50'b11_1011110000010111_0111110000010011_1111110000010111;
      patterns[2900] = 50'b00_1100100001111101_0101101100000010_0010001101111111;
      patterns[2901] = 50'b01_1100100001111101_0101101100000010_0110110101111011;
      patterns[2902] = 50'b10_1100100001111101_0101101100000010_0100100000000000;
      patterns[2903] = 50'b11_1100100001111101_0101101100000010_1101101101111111;
      patterns[2904] = 50'b00_1101101111001000_0010100101100110_0000010100101110;
      patterns[2905] = 50'b01_1101101111001000_0010100101100110_1011001001100010;
      patterns[2906] = 50'b10_1101101111001000_0010100101100110_0000100101000000;
      patterns[2907] = 50'b11_1101101111001000_0010100101100110_1111101111101110;
      patterns[2908] = 50'b00_0101100111101111_0100000001100111_1001101001010110;
      patterns[2909] = 50'b01_0101100111101111_0100000001100111_0001100110001000;
      patterns[2910] = 50'b10_0101100111101111_0100000001100111_0100000001100111;
      patterns[2911] = 50'b11_0101100111101111_0100000001100111_0101100111101111;
      patterns[2912] = 50'b00_0111011101000100_1010111101011001_0010011010011101;
      patterns[2913] = 50'b01_0111011101000100_1010111101011001_1100011111101011;
      patterns[2914] = 50'b10_0111011101000100_1010111101011001_0010011101000000;
      patterns[2915] = 50'b11_0111011101000100_1010111101011001_1111111101011101;
      patterns[2916] = 50'b00_1100100111000111_0010000010100001_1110101001101000;
      patterns[2917] = 50'b01_1100100111000111_0010000010100001_1010100100100110;
      patterns[2918] = 50'b10_1100100111000111_0010000010100001_0000000010000001;
      patterns[2919] = 50'b11_1100100111000111_0010000010100001_1110100111100111;
      patterns[2920] = 50'b00_0000000110110000_1100111010001111_1101000000111111;
      patterns[2921] = 50'b01_0000000110110000_1100111010001111_0011001100100001;
      patterns[2922] = 50'b10_0000000110110000_1100111010001111_0000000010000000;
      patterns[2923] = 50'b11_0000000110110000_1100111010001111_1100111110111111;
      patterns[2924] = 50'b00_1100011111000001_1000111100000100_0101011011000101;
      patterns[2925] = 50'b01_1100011111000001_1000111100000100_0011100010111101;
      patterns[2926] = 50'b10_1100011111000001_1000111100000100_1000011100000000;
      patterns[2927] = 50'b11_1100011111000001_1000111100000100_1100111111000101;
      patterns[2928] = 50'b00_0000010100111001_0010000010111101_0010010111110110;
      patterns[2929] = 50'b01_0000010100111001_0010000010111101_1110010001111100;
      patterns[2930] = 50'b10_0000010100111001_0010000010111101_0000000000111001;
      patterns[2931] = 50'b11_0000010100111001_0010000010111101_0010010110111101;
      patterns[2932] = 50'b00_0011101111100101_1111001011100011_0010111011001000;
      patterns[2933] = 50'b01_0011101111100101_1111001011100011_0100100100000010;
      patterns[2934] = 50'b10_0011101111100101_1111001011100011_0011001011100001;
      patterns[2935] = 50'b11_0011101111100101_1111001011100011_1111101111100111;
      patterns[2936] = 50'b00_1101101001111010_1111111000101110_1101100010101000;
      patterns[2937] = 50'b01_1101101001111010_1111111000101110_1101110001001100;
      patterns[2938] = 50'b10_1101101001111010_1111111000101110_1101101000101010;
      patterns[2939] = 50'b11_1101101001111010_1111111000101110_1111111001111110;
      patterns[2940] = 50'b00_0111101011110100_1001000111101000_0000110011011100;
      patterns[2941] = 50'b01_0111101011110100_1001000111101000_1110100100001100;
      patterns[2942] = 50'b10_0111101011110100_1001000111101000_0001000011100000;
      patterns[2943] = 50'b11_0111101011110100_1001000111101000_1111101111111100;
      patterns[2944] = 50'b00_1110001111001110_0011110101100110_0010000100110100;
      patterns[2945] = 50'b01_1110001111001110_0011110101100110_1010011001101000;
      patterns[2946] = 50'b10_1110001111001110_0011110101100110_0010000101000110;
      patterns[2947] = 50'b11_1110001111001110_0011110101100110_1111111111101110;
      patterns[2948] = 50'b00_0011101001100100_0000001110110111_0011111000011011;
      patterns[2949] = 50'b01_0011101001100100_0000001110110111_0011011010101101;
      patterns[2950] = 50'b10_0011101001100100_0000001110110111_0000001000100100;
      patterns[2951] = 50'b11_0011101001100100_0000001110110111_0011101111110111;
      patterns[2952] = 50'b00_1010101000110111_1000001000110010_0010110001101001;
      patterns[2953] = 50'b01_1010101000110111_1000001000110010_0010100000000101;
      patterns[2954] = 50'b10_1010101000110111_1000001000110010_1000001000110010;
      patterns[2955] = 50'b11_1010101000110111_1000001000110010_1010101000110111;
      patterns[2956] = 50'b00_1000001101010011_1000111011101011_0001001000111110;
      patterns[2957] = 50'b01_1000001101010011_1000111011101011_1111010001101000;
      patterns[2958] = 50'b10_1000001101010011_1000111011101011_1000001001000011;
      patterns[2959] = 50'b11_1000001101010011_1000111011101011_1000111111111011;
      patterns[2960] = 50'b00_0111011011010101_0111000010101010_1110011101111111;
      patterns[2961] = 50'b01_0111011011010101_0111000010101010_0000011000101011;
      patterns[2962] = 50'b10_0111011011010101_0111000010101010_0111000010000000;
      patterns[2963] = 50'b11_0111011011010101_0111000010101010_0111011011111111;
      patterns[2964] = 50'b00_1011010011110110_0100001001110011_1111011101101001;
      patterns[2965] = 50'b01_1011010011110110_0100001001110011_0111001010000011;
      patterns[2966] = 50'b10_1011010011110110_0100001001110011_0000000001110010;
      patterns[2967] = 50'b11_1011010011110110_0100001001110011_1111011011110111;
      patterns[2968] = 50'b00_1010100100110010_0101111111110110_0000100100101000;
      patterns[2969] = 50'b01_1010100100110010_0101111111110110_0100100100111100;
      patterns[2970] = 50'b10_1010100100110010_0101111111110110_0000100100110010;
      patterns[2971] = 50'b11_1010100100110010_0101111111110110_1111111111110110;
      patterns[2972] = 50'b00_0110000001111001_0001100111011101_0111101001010110;
      patterns[2973] = 50'b01_0110000001111001_0001100111011101_0100011010011100;
      patterns[2974] = 50'b10_0110000001111001_0001100111011101_0000000001011001;
      patterns[2975] = 50'b11_0110000001111001_0001100111011101_0111100111111101;
      patterns[2976] = 50'b00_0001011111010101_0001011111011010_0010111110101111;
      patterns[2977] = 50'b01_0001011111010101_0001011111011010_1111111111111011;
      patterns[2978] = 50'b10_0001011111010101_0001011111011010_0001011111010000;
      patterns[2979] = 50'b11_0001011111010101_0001011111011010_0001011111011111;
      patterns[2980] = 50'b00_0110100101010101_0001111000010111_1000011101101100;
      patterns[2981] = 50'b01_0110100101010101_0001111000010111_0100101100111110;
      patterns[2982] = 50'b10_0110100101010101_0001111000010111_0000100000010101;
      patterns[2983] = 50'b11_0110100101010101_0001111000010111_0111111101010111;
      patterns[2984] = 50'b00_0011110111010100_1011101101001110_1111100100100010;
      patterns[2985] = 50'b01_0011110111010100_1011101101001110_1000001010000110;
      patterns[2986] = 50'b10_0011110111010100_1011101101001110_0011100101000100;
      patterns[2987] = 50'b11_0011110111010100_1011101101001110_1011111111011110;
      patterns[2988] = 50'b00_0101111010000010_0011111110100111_1001111000101001;
      patterns[2989] = 50'b01_0101111010000010_0011111110100111_0001111011011011;
      patterns[2990] = 50'b10_0101111010000010_0011111110100111_0001111010000010;
      patterns[2991] = 50'b11_0101111010000010_0011111110100111_0111111110100111;
      patterns[2992] = 50'b00_1101010101100100_0100000111000011_0001011100100111;
      patterns[2993] = 50'b01_1101010101100100_0100000111000011_1001001110100001;
      patterns[2994] = 50'b10_1101010101100100_0100000111000011_0100000101000000;
      patterns[2995] = 50'b11_1101010101100100_0100000111000011_1101010111100111;
      patterns[2996] = 50'b00_0111001000001111_1001101001111111_0000110010001110;
      patterns[2997] = 50'b01_0111001000001111_1001101001111111_1101011110010000;
      patterns[2998] = 50'b10_0111001000001111_1001101001111111_0001001000001111;
      patterns[2999] = 50'b11_0111001000001111_1001101001111111_1111101001111111;
      patterns[3000] = 50'b00_1100010010100011_1100011110111100_1000110001011111;
      patterns[3001] = 50'b01_1100010010100011_1100011110111100_1111110011100111;
      patterns[3002] = 50'b10_1100010010100011_1100011110111100_1100010010100000;
      patterns[3003] = 50'b11_1100010010100011_1100011110111100_1100011110111111;
      patterns[3004] = 50'b00_1100111000011000_1110111011010010_1011110011101010;
      patterns[3005] = 50'b01_1100111000011000_1110111011010010_1101111101000110;
      patterns[3006] = 50'b10_1100111000011000_1110111011010010_1100111000010000;
      patterns[3007] = 50'b11_1100111000011000_1110111011010010_1110111011011010;
      patterns[3008] = 50'b00_1110111100001010_1000111011100100_0111110111101110;
      patterns[3009] = 50'b01_1110111100001010_1000111011100100_0110000000100110;
      patterns[3010] = 50'b10_1110111100001010_1000111011100100_1000111000000000;
      patterns[3011] = 50'b11_1110111100001010_1000111011100100_1110111111101110;
      patterns[3012] = 50'b00_0100011100010000_0101110110010011_1010010010100011;
      patterns[3013] = 50'b01_0100011100010000_0101110110010011_1110100101111101;
      patterns[3014] = 50'b10_0100011100010000_0101110110010011_0100010100010000;
      patterns[3015] = 50'b11_0100011100010000_0101110110010011_0101111110010011;
      patterns[3016] = 50'b00_1001001101010100_1011110011011111_0101000000110011;
      patterns[3017] = 50'b01_1001001101010100_1011110011011111_1101011001110101;
      patterns[3018] = 50'b10_1001001101010100_1011110011011111_1001000001010100;
      patterns[3019] = 50'b11_1001001101010100_1011110011011111_1011111111011111;
      patterns[3020] = 50'b00_1001010011010100_1110001010010010_0111011101100110;
      patterns[3021] = 50'b01_1001010011010100_1110001010010010_1011001001000010;
      patterns[3022] = 50'b10_1001010011010100_1110001010010010_1000000010010000;
      patterns[3023] = 50'b11_1001010011010100_1110001010010010_1111011011010110;
      patterns[3024] = 50'b00_0101101010111111_1100011101010100_0010001000010011;
      patterns[3025] = 50'b01_0101101010111111_1100011101010100_1001001101101011;
      patterns[3026] = 50'b10_0101101010111111_1100011101010100_0100001000010100;
      patterns[3027] = 50'b11_0101101010111111_1100011101010100_1101111111111111;
      patterns[3028] = 50'b00_0100110100010010_1001100101011010_1110011001101100;
      patterns[3029] = 50'b01_0100110100010010_1001100101011010_1011001110111000;
      patterns[3030] = 50'b10_0100110100010010_1001100101011010_0000100100010010;
      patterns[3031] = 50'b11_0100110100010010_1001100101011010_1101110101011010;
      patterns[3032] = 50'b00_0010001111110010_0000001100011000_0010011100001010;
      patterns[3033] = 50'b01_0010001111110010_0000001100011000_0010000011011010;
      patterns[3034] = 50'b10_0010001111110010_0000001100011000_0000001100010000;
      patterns[3035] = 50'b11_0010001111110010_0000001100011000_0010001111111010;
      patterns[3036] = 50'b00_1101001011101011_1001010100111000_0110100000100011;
      patterns[3037] = 50'b01_1101001011101011_1001010100111000_0011110110110011;
      patterns[3038] = 50'b10_1101001011101011_1001010100111000_1001000000101000;
      patterns[3039] = 50'b11_1101001011101011_1001010100111000_1101011111111011;
      patterns[3040] = 50'b00_1110000011111011_1111101101011110_1101110001011001;
      patterns[3041] = 50'b01_1110000011111011_1111101101011110_1110010110011101;
      patterns[3042] = 50'b10_1110000011111011_1111101101011110_1110000001011010;
      patterns[3043] = 50'b11_1110000011111011_1111101101011110_1111101111111111;
      patterns[3044] = 50'b00_0101000011010111_1111100000010111_0100100011101110;
      patterns[3045] = 50'b01_0101000011010111_1111100000010111_0101100011000000;
      patterns[3046] = 50'b10_0101000011010111_1111100000010111_0101000000010111;
      patterns[3047] = 50'b11_0101000011010111_1111100000010111_1111100011010111;
      patterns[3048] = 50'b00_1001010100010111_0000110101011110_1010001001110101;
      patterns[3049] = 50'b01_1001010100010111_0000110101011110_1000011110111001;
      patterns[3050] = 50'b10_1001010100010111_0000110101011110_0000010100010110;
      patterns[3051] = 50'b11_1001010100010111_0000110101011110_1001110101011111;
      patterns[3052] = 50'b00_1001101100111100_1111111100100001_1001101001011101;
      patterns[3053] = 50'b01_1001101100111100_1111111100100001_1001110000011011;
      patterns[3054] = 50'b10_1001101100111100_1111111100100001_1001101100100000;
      patterns[3055] = 50'b11_1001101100111100_1111111100100001_1111111100111101;
      patterns[3056] = 50'b00_1001110001010111_0100001111010100_1110000000101011;
      patterns[3057] = 50'b01_1001110001010111_0100001111010100_0101100010000011;
      patterns[3058] = 50'b10_1001110001010111_0100001111010100_0000000001010100;
      patterns[3059] = 50'b11_1001110001010111_0100001111010100_1101111111010111;
      patterns[3060] = 50'b00_1000101100111011_1110111101000101_0111101010000000;
      patterns[3061] = 50'b01_1000101100111011_1110111101000101_1001101111110110;
      patterns[3062] = 50'b10_1000101100111011_1110111101000101_1000101100000001;
      patterns[3063] = 50'b11_1000101100111011_1110111101000101_1110111101111111;
      patterns[3064] = 50'b00_1110110000111000_1001010101001001_1000000110000001;
      patterns[3065] = 50'b01_1110110000111000_1001010101001001_0101011011101111;
      patterns[3066] = 50'b10_1110110000111000_1001010101001001_1000010000001000;
      patterns[3067] = 50'b11_1110110000111000_1001010101001001_1111110101111001;
      patterns[3068] = 50'b00_1111101010100100_0010011100010011_0010000110110111;
      patterns[3069] = 50'b01_1111101010100100_0010011100010011_1101001110010001;
      patterns[3070] = 50'b10_1111101010100100_0010011100010011_0010001000000000;
      patterns[3071] = 50'b11_1111101010100100_0010011100010011_1111111110110111;
      patterns[3072] = 50'b00_1110100111001010_0111011100010000_0110000011011010;
      patterns[3073] = 50'b01_1110100111001010_0111011100010000_0111001010111010;
      patterns[3074] = 50'b10_1110100111001010_0111011100010000_0110000100000000;
      patterns[3075] = 50'b11_1110100111001010_0111011100010000_1111111111011010;
      patterns[3076] = 50'b00_0000101100010110_0001111010010101_0010100110101011;
      patterns[3077] = 50'b01_0000101100010110_0001111010010101_1110110010000001;
      patterns[3078] = 50'b10_0000101100010110_0001111010010101_0000101000010100;
      patterns[3079] = 50'b11_0000101100010110_0001111010010101_0001111110010111;
      patterns[3080] = 50'b00_1100011100001010_0010111001010001_1111010101011011;
      patterns[3081] = 50'b01_1100011100001010_0010111001010001_1001100010111001;
      patterns[3082] = 50'b10_1100011100001010_0010111001010001_0000011000000000;
      patterns[3083] = 50'b11_1100011100001010_0010111001010001_1110111101011011;
      patterns[3084] = 50'b00_1100101110110010_1100100100010001_1001010011000011;
      patterns[3085] = 50'b01_1100101110110010_1100100100010001_0000001010100001;
      patterns[3086] = 50'b10_1100101110110010_1100100100010001_1100100100010000;
      patterns[3087] = 50'b11_1100101110110010_1100100100010001_1100101110110011;
      patterns[3088] = 50'b00_0001011001110001_0110011110101110_0111111000011111;
      patterns[3089] = 50'b01_0001011001110001_0110011110101110_1010111011000011;
      patterns[3090] = 50'b10_0001011001110001_0110011110101110_0000011000100000;
      patterns[3091] = 50'b11_0001011001110001_0110011110101110_0111011111111111;
      patterns[3092] = 50'b00_1010000111111001_1001111111011010_0100000111010011;
      patterns[3093] = 50'b01_1010000111111001_1001111111011010_0000001000011111;
      patterns[3094] = 50'b10_1010000111111001_1001111111011010_1000000111011000;
      patterns[3095] = 50'b11_1010000111111001_1001111111011010_1011111111111011;
      patterns[3096] = 50'b00_0110100011110101_0110010100111111_1100111000110100;
      patterns[3097] = 50'b01_0110100011110101_0110010100111111_0000001110110110;
      patterns[3098] = 50'b10_0110100011110101_0110010100111111_0110000000110101;
      patterns[3099] = 50'b11_0110100011110101_0110010100111111_0110110111111111;
      patterns[3100] = 50'b00_0001001110101000_1001100010100001_1010110001001001;
      patterns[3101] = 50'b01_0001001110101000_1001100010100001_0111101100000111;
      patterns[3102] = 50'b10_0001001110101000_1001100010100001_0001000010100000;
      patterns[3103] = 50'b11_0001001110101000_1001100010100001_1001101110101001;
      patterns[3104] = 50'b00_0101011111101110_1000000111111011_1101100111101001;
      patterns[3105] = 50'b01_0101011111101110_1000000111111011_1101010111110011;
      patterns[3106] = 50'b10_0101011111101110_1000000111111011_0000000111101010;
      patterns[3107] = 50'b11_0101011111101110_1000000111111011_1101011111111111;
      patterns[3108] = 50'b00_1011000010111000_0110110011101010_0001110110100010;
      patterns[3109] = 50'b01_1011000010111000_0110110011101010_0100001111001110;
      patterns[3110] = 50'b10_1011000010111000_0110110011101010_0010000010101000;
      patterns[3111] = 50'b11_1011000010111000_0110110011101010_1111110011111010;
      patterns[3112] = 50'b00_0101000110100000_1110000011010100_0011001001110100;
      patterns[3113] = 50'b01_0101000110100000_1110000011010100_0111000011001100;
      patterns[3114] = 50'b10_0101000110100000_1110000011010100_0100000010000000;
      patterns[3115] = 50'b11_0101000110100000_1110000011010100_1111000111110100;
      patterns[3116] = 50'b00_1110010111010000_1110001110001100_1100100101011100;
      patterns[3117] = 50'b01_1110010111010000_1110001110001100_0000001001000100;
      patterns[3118] = 50'b10_1110010111010000_1110001110001100_1110000110000000;
      patterns[3119] = 50'b11_1110010111010000_1110001110001100_1110011111011100;
      patterns[3120] = 50'b00_1101110001011111_1101110100001111_1011100101101110;
      patterns[3121] = 50'b01_1101110001011111_1101110100001111_1111111101010000;
      patterns[3122] = 50'b10_1101110001011111_1101110100001111_1101110000001111;
      patterns[3123] = 50'b11_1101110001011111_1101110100001111_1101110101011111;
      patterns[3124] = 50'b00_0111000011001011_0100000001110101_1011000101000000;
      patterns[3125] = 50'b01_0111000011001011_0100000001110101_0011000001010110;
      patterns[3126] = 50'b10_0111000011001011_0100000001110101_0100000001000001;
      patterns[3127] = 50'b11_0111000011001011_0100000001110101_0111000011111111;
      patterns[3128] = 50'b00_1100100110001101_0011100010100011_0000001000110000;
      patterns[3129] = 50'b01_1100100110001101_0011100010100011_1001000011101010;
      patterns[3130] = 50'b10_1100100110001101_0011100010100011_0000100010000001;
      patterns[3131] = 50'b11_1100100110001101_0011100010100011_1111100110101111;
      patterns[3132] = 50'b00_0000101000101010_1001101000000111_1010010000110001;
      patterns[3133] = 50'b01_0000101000101010_1001101000000111_0111000000100011;
      patterns[3134] = 50'b10_0000101000101010_1001101000000111_0000101000000010;
      patterns[3135] = 50'b11_0000101000101010_1001101000000111_1001101000101111;
      patterns[3136] = 50'b00_1111111011100100_0001010010100111_0001001110001011;
      patterns[3137] = 50'b01_1111111011100100_0001010010100111_1110101000111101;
      patterns[3138] = 50'b10_1111111011100100_0001010010100111_0001010010100100;
      patterns[3139] = 50'b11_1111111011100100_0001010010100111_1111111011100111;
      patterns[3140] = 50'b00_1001011110000101_1001011011001011_0010111001010000;
      patterns[3141] = 50'b01_1001011110000101_1001011011001011_0000000010111010;
      patterns[3142] = 50'b10_1001011110000101_1001011011001011_1001011010000001;
      patterns[3143] = 50'b11_1001011110000101_1001011011001011_1001011111001111;
      patterns[3144] = 50'b00_0001000111001101_0111011100100000_1000100011101101;
      patterns[3145] = 50'b01_0001000111001101_0111011100100000_1001101010101101;
      patterns[3146] = 50'b10_0001000111001101_0111011100100000_0001000100000000;
      patterns[3147] = 50'b11_0001000111001101_0111011100100000_0111011111101101;
      patterns[3148] = 50'b00_1110010001100111_0000000101011001_1110010111000000;
      patterns[3149] = 50'b01_1110010001100111_0000000101011001_1110001100001110;
      patterns[3150] = 50'b10_1110010001100111_0000000101011001_0000000001000001;
      patterns[3151] = 50'b11_1110010001100111_0000000101011001_1110010101111111;
      patterns[3152] = 50'b00_1110110110111011_1000000010101011_0110111001100110;
      patterns[3153] = 50'b01_1110110110111011_1000000010101011_0110110100010000;
      patterns[3154] = 50'b10_1110110110111011_1000000010101011_1000000010101011;
      patterns[3155] = 50'b11_1110110110111011_1000000010101011_1110110110111011;
      patterns[3156] = 50'b00_0111000000011001_1011001110011111_0010001110111000;
      patterns[3157] = 50'b01_0111000000011001_1011001110011111_1011110001111010;
      patterns[3158] = 50'b10_0111000000011001_1011001110011111_0011000000011001;
      patterns[3159] = 50'b11_0111000000011001_1011001110011111_1111001110011111;
      patterns[3160] = 50'b00_0010001111000011_0111101111100010_1001111110100101;
      patterns[3161] = 50'b01_0010001111000011_0111101111100010_1010011111100001;
      patterns[3162] = 50'b10_0010001111000011_0111101111100010_0010001111000010;
      patterns[3163] = 50'b11_0010001111000011_0111101111100010_0111101111100011;
      patterns[3164] = 50'b00_0101100001000010_1001010111110110_1110111000111000;
      patterns[3165] = 50'b01_0101100001000010_1001010111110110_1100001001001100;
      patterns[3166] = 50'b10_0101100001000010_1001010111110110_0001000001000010;
      patterns[3167] = 50'b11_0101100001000010_1001010111110110_1101110111110110;
      patterns[3168] = 50'b00_0100111011110000_1001111101101011_1110111001011011;
      patterns[3169] = 50'b01_0100111011110000_1001111101101011_1010111110000101;
      patterns[3170] = 50'b10_0100111011110000_1001111101101011_0000111001100000;
      patterns[3171] = 50'b11_0100111011110000_1001111101101011_1101111111111011;
      patterns[3172] = 50'b00_1100100101111011_1101000110110001_1001101100101100;
      patterns[3173] = 50'b01_1100100101111011_1101000110110001_1111011111001010;
      patterns[3174] = 50'b10_1100100101111011_1101000110110001_1100000100110001;
      patterns[3175] = 50'b11_1100100101111011_1101000110110001_1101100111111011;
      patterns[3176] = 50'b00_0010111000000001_1011001100011000_1110000100011001;
      patterns[3177] = 50'b01_0010111000000001_1011001100011000_0111101011101001;
      patterns[3178] = 50'b10_0010111000000001_1011001100011000_0010001000000000;
      patterns[3179] = 50'b11_0010111000000001_1011001100011000_1011111100011001;
      patterns[3180] = 50'b00_1010100000100000_1110001000000011_1000101000100011;
      patterns[3181] = 50'b01_1010100000100000_1110001000000011_1100011000011101;
      patterns[3182] = 50'b10_1010100000100000_1110001000000011_1010000000000000;
      patterns[3183] = 50'b11_1010100000100000_1110001000000011_1110101000100011;
      patterns[3184] = 50'b00_1011000010100000_1100011110001100_0111100000101100;
      patterns[3185] = 50'b01_1011000010100000_1100011110001100_1110100100010100;
      patterns[3186] = 50'b10_1011000010100000_1100011110001100_1000000010000000;
      patterns[3187] = 50'b11_1011000010100000_1100011110001100_1111011110101100;
      patterns[3188] = 50'b00_0101010100001100_1110000101111001_0011011010000101;
      patterns[3189] = 50'b01_0101010100001100_1110000101111001_0111001110010011;
      patterns[3190] = 50'b10_0101010100001100_1110000101111001_0100000100001000;
      patterns[3191] = 50'b11_0101010100001100_1110000101111001_1111010101111101;
      patterns[3192] = 50'b00_0011101100110010_1101011100110110_0001001001101000;
      patterns[3193] = 50'b01_0011101100110010_1101011100110110_0110001111111100;
      patterns[3194] = 50'b10_0011101100110010_1101011100110110_0001001100110010;
      patterns[3195] = 50'b11_0011101100110010_1101011100110110_1111111100110110;
      patterns[3196] = 50'b00_1000101100001101_0100110101011100_1101100001101001;
      patterns[3197] = 50'b01_1000101100001101_0100110101011100_0011110110110001;
      patterns[3198] = 50'b10_1000101100001101_0100110101011100_0000100100001100;
      patterns[3199] = 50'b11_1000101100001101_0100110101011100_1100111101011101;
      patterns[3200] = 50'b00_1101000111010010_0111011010110011_0100100010000101;
      patterns[3201] = 50'b01_1101000111010010_0111011010110011_0101101100011111;
      patterns[3202] = 50'b10_1101000111010010_0111011010110011_0101000010010010;
      patterns[3203] = 50'b11_1101000111010010_0111011010110011_1111011111110011;
      patterns[3204] = 50'b00_0101001100100110_0111101110111110_1100111011100100;
      patterns[3205] = 50'b01_0101001100100110_0111101110111110_1101011101101000;
      patterns[3206] = 50'b10_0101001100100110_0111101110111110_0101001100100110;
      patterns[3207] = 50'b11_0101001100100110_0111101110111110_0111101110111110;
      patterns[3208] = 50'b00_1011000000011111_1011000111010010_0110000111110001;
      patterns[3209] = 50'b01_1011000000011111_1011000111010010_1111111001001101;
      patterns[3210] = 50'b10_1011000000011111_1011000111010010_1011000000010010;
      patterns[3211] = 50'b11_1011000000011111_1011000111010010_1011000111011111;
      patterns[3212] = 50'b00_1111011100001110_0010110000000010_0010001100010000;
      patterns[3213] = 50'b01_1111011100001110_0010110000000010_1100101100001100;
      patterns[3214] = 50'b10_1111011100001110_0010110000000010_0010010000000010;
      patterns[3215] = 50'b11_1111011100001110_0010110000000010_1111111100001110;
      patterns[3216] = 50'b00_0001000011100011_1101000111010111_1110001010111010;
      patterns[3217] = 50'b01_0001000011100011_1101000111010111_0011111100001100;
      patterns[3218] = 50'b10_0001000011100011_1101000111010111_0001000011000011;
      patterns[3219] = 50'b11_0001000011100011_1101000111010111_1101000111110111;
      patterns[3220] = 50'b00_1010101001101100_1110110100100011_1001011110001111;
      patterns[3221] = 50'b01_1010101001101100_1110110100100011_1011110101001001;
      patterns[3222] = 50'b10_1010101001101100_1110110100100011_1010100000100000;
      patterns[3223] = 50'b11_1010101001101100_1110110100100011_1110111101101111;
      patterns[3224] = 50'b00_1000110111000101_0001000010110100_1001111001111001;
      patterns[3225] = 50'b01_1000110111000101_0001000010110100_0111110100010001;
      patterns[3226] = 50'b10_1000110111000101_0001000010110100_0000000010000100;
      patterns[3227] = 50'b11_1000110111000101_0001000010110100_1001110111110101;
      patterns[3228] = 50'b00_0101110010111111_1001000000001000_1110110011000111;
      patterns[3229] = 50'b01_0101110010111111_1001000000001000_1100110010110111;
      patterns[3230] = 50'b10_0101110010111111_1001000000001000_0001000000001000;
      patterns[3231] = 50'b11_0101110010111111_1001000000001000_1101110010111111;
      patterns[3232] = 50'b00_1000110010000101_0010110001010000_1011100011010101;
      patterns[3233] = 50'b01_1000110010000101_0010110001010000_0110000000110101;
      patterns[3234] = 50'b10_1000110010000101_0010110001010000_0000110000000000;
      patterns[3235] = 50'b11_1000110010000101_0010110001010000_1010110011010101;
      patterns[3236] = 50'b00_1100011011111101_0111111110101010_0100011010100111;
      patterns[3237] = 50'b01_1100011011111101_0111111110101010_0100011101010011;
      patterns[3238] = 50'b10_1100011011111101_0111111110101010_0100011010101000;
      patterns[3239] = 50'b11_1100011011111101_0111111110101010_1111111111111111;
      patterns[3240] = 50'b00_1010010001111011_0110010000100000_0000100010011011;
      patterns[3241] = 50'b01_1010010001111011_0110010000100000_0100000001011011;
      patterns[3242] = 50'b10_1010010001111011_0110010000100000_0010010000100000;
      patterns[3243] = 50'b11_1010010001111011_0110010000100000_1110010001111011;
      patterns[3244] = 50'b00_0101000101001110_1010001111100111_1111010100110101;
      patterns[3245] = 50'b01_0101000101001110_1010001111100111_1010110101100111;
      patterns[3246] = 50'b10_0101000101001110_1010001111100111_0000000101000110;
      patterns[3247] = 50'b11_0101000101001110_1010001111100111_1111001111101111;
      patterns[3248] = 50'b00_1100010001010001_1010101010011001_0110111011101010;
      patterns[3249] = 50'b01_1100010001010001_1010101010011001_0001100110111000;
      patterns[3250] = 50'b10_1100010001010001_1010101010011001_1000000000010001;
      patterns[3251] = 50'b11_1100010001010001_1010101010011001_1110111011011001;
      patterns[3252] = 50'b00_1101111001110100_0110011100101000_0100010110011100;
      patterns[3253] = 50'b01_1101111001110100_0110011100101000_0111011101001100;
      patterns[3254] = 50'b10_1101111001110100_0110011100101000_0100011000100000;
      patterns[3255] = 50'b11_1101111001110100_0110011100101000_1111111101111100;
      patterns[3256] = 50'b00_0010010100110100_1011101101001111_1110000010000011;
      patterns[3257] = 50'b01_0010010100110100_1011101101001111_0110100111100101;
      patterns[3258] = 50'b10_0010010100110100_1011101101001111_0010000100000100;
      patterns[3259] = 50'b11_0010010100110100_1011101101001111_1011111101111111;
      patterns[3260] = 50'b00_1110001111000011_1001001001010101_0111011000011000;
      patterns[3261] = 50'b01_1110001111000011_1001001001010101_0101000101101110;
      patterns[3262] = 50'b10_1110001111000011_1001001001010101_1000001001000001;
      patterns[3263] = 50'b11_1110001111000011_1001001001010101_1111001111010111;
      patterns[3264] = 50'b00_1100010111110100_0101010111000000_0001101110110100;
      patterns[3265] = 50'b01_1100010111110100_0101010111000000_0111000000110100;
      patterns[3266] = 50'b10_1100010111110100_0101010111000000_0100010111000000;
      patterns[3267] = 50'b11_1100010111110100_0101010111000000_1101010111110100;
      patterns[3268] = 50'b00_0111010110111010_1111010110101111_0110101101101001;
      patterns[3269] = 50'b01_0111010110111010_1111010110101111_1000000000001011;
      patterns[3270] = 50'b10_0111010110111010_1111010110101111_0111010110101010;
      patterns[3271] = 50'b11_0111010110111010_1111010110101111_1111010110111111;
      patterns[3272] = 50'b00_0011110111001111_0001010000011100_0101000111101011;
      patterns[3273] = 50'b01_0011110111001111_0001010000011100_0010100110110011;
      patterns[3274] = 50'b10_0011110111001111_0001010000011100_0001010000001100;
      patterns[3275] = 50'b11_0011110111001111_0001010000011100_0011110111011111;
      patterns[3276] = 50'b00_0001101010100000_0100000010000100_0101101100100100;
      patterns[3277] = 50'b01_0001101010100000_0100000010000100_1101101000011100;
      patterns[3278] = 50'b10_0001101010100000_0100000010000100_0000000010000000;
      patterns[3279] = 50'b11_0001101010100000_0100000010000100_0101101010100100;
      patterns[3280] = 50'b00_0011001111100100_0011010010010010_0110100001110110;
      patterns[3281] = 50'b01_0011001111100100_0011010010010010_1111111101010010;
      patterns[3282] = 50'b10_0011001111100100_0011010010010010_0011000010000000;
      patterns[3283] = 50'b11_0011001111100100_0011010010010010_0011011111110110;
      patterns[3284] = 50'b00_0100010110110011_1111110011101001_0100001010011100;
      patterns[3285] = 50'b01_0100010110110011_1111110011101001_0100100011001010;
      patterns[3286] = 50'b10_0100010110110011_1111110011101001_0100010010100001;
      patterns[3287] = 50'b11_0100010110110011_1111110011101001_1111110111111011;
      patterns[3288] = 50'b00_1010110101111101_0011001011101000_1110000001100101;
      patterns[3289] = 50'b01_1010110101111101_0011001011101000_0111101010010101;
      patterns[3290] = 50'b10_1010110101111101_0011001011101000_0010000001101000;
      patterns[3291] = 50'b11_1010110101111101_0011001011101000_1011111111111101;
      patterns[3292] = 50'b00_0101011011010011_0101111111011001_1011011010101100;
      patterns[3293] = 50'b01_0101011011010011_0101111111011001_1111011011111010;
      patterns[3294] = 50'b10_0101011011010011_0101111111011001_0101011011010001;
      patterns[3295] = 50'b11_0101011011010011_0101111111011001_0101111111011011;
      patterns[3296] = 50'b00_1011001010110111_0011111101110101_1111001000101100;
      patterns[3297] = 50'b01_1011001010110111_0011111101110101_0111001101000010;
      patterns[3298] = 50'b10_1011001010110111_0011111101110101_0011001000110101;
      patterns[3299] = 50'b11_1011001010110111_0011111101110101_1011111111110111;
      patterns[3300] = 50'b00_1101101110110110_1000000101101110_0101110100100100;
      patterns[3301] = 50'b01_1101101110110110_1000000101101110_0101101001001000;
      patterns[3302] = 50'b10_1101101110110110_1000000101101110_1000000100100110;
      patterns[3303] = 50'b11_1101101110110110_1000000101101110_1101101111111110;
      patterns[3304] = 50'b00_0111111000111011_0111011110110001_1111010111101100;
      patterns[3305] = 50'b01_0111111000111011_0111011110110001_0000011010001010;
      patterns[3306] = 50'b10_0111111000111011_0111011110110001_0111011000110001;
      patterns[3307] = 50'b11_0111111000111011_0111011110110001_0111111110111011;
      patterns[3308] = 50'b00_1001100011111111_1001110000011001_0011010100011000;
      patterns[3309] = 50'b01_1001100011111111_1001110000011001_1111110011100110;
      patterns[3310] = 50'b10_1001100011111111_1001110000011001_1001100000011001;
      patterns[3311] = 50'b11_1001100011111111_1001110000011001_1001110011111111;
      patterns[3312] = 50'b00_1000101000000001_0100001111111011_1100110111111100;
      patterns[3313] = 50'b01_1000101000000001_0100001111111011_0100011000000110;
      patterns[3314] = 50'b10_1000101000000001_0100001111111011_0000001000000001;
      patterns[3315] = 50'b11_1000101000000001_0100001111111011_1100101111111011;
      patterns[3316] = 50'b00_1001001011100001_0010010100000101_1011011111100110;
      patterns[3317] = 50'b01_1001001011100001_0010010100000101_0110110111011100;
      patterns[3318] = 50'b10_1001001011100001_0010010100000101_0000000000000001;
      patterns[3319] = 50'b11_1001001011100001_0010010100000101_1011011111100101;
      patterns[3320] = 50'b00_0101000001011110_0110010101010111_1011010110110101;
      patterns[3321] = 50'b01_0101000001011110_0110010101010111_1110101100000111;
      patterns[3322] = 50'b10_0101000001011110_0110010101010111_0100000001010110;
      patterns[3323] = 50'b11_0101000001011110_0110010101010111_0111010101011111;
      patterns[3324] = 50'b00_1110011000010010_1110101100001000_1101000100011010;
      patterns[3325] = 50'b01_1110011000010010_1110101100001000_1111101100001010;
      patterns[3326] = 50'b10_1110011000010010_1110101100001000_1110001000000000;
      patterns[3327] = 50'b11_1110011000010010_1110101100001000_1110111100011010;
      patterns[3328] = 50'b00_1000010111001110_0000110100100100_1001001011110010;
      patterns[3329] = 50'b01_1000010111001110_0000110100100100_0111100010101010;
      patterns[3330] = 50'b10_1000010111001110_0000110100100100_0000010100000100;
      patterns[3331] = 50'b11_1000010111001110_0000110100100100_1000110111101110;
      patterns[3332] = 50'b00_1100001100111110_1110110011011110_1011000000011100;
      patterns[3333] = 50'b01_1100001100111110_1110110011011110_1101011001100000;
      patterns[3334] = 50'b10_1100001100111110_1110110011011110_1100000000011110;
      patterns[3335] = 50'b11_1100001100111110_1110110011011110_1110111111111110;
      patterns[3336] = 50'b00_1110010100111001_1101000000100011_1011010101011100;
      patterns[3337] = 50'b01_1110010100111001_1101000000100011_0001010100010110;
      patterns[3338] = 50'b10_1110010100111001_1101000000100011_1100000000100001;
      patterns[3339] = 50'b11_1110010100111001_1101000000100011_1111010100111011;
      patterns[3340] = 50'b00_0100100000111011_0100001001111100_1000101010110111;
      patterns[3341] = 50'b01_0100100000111011_0100001001111100_0000010110111111;
      patterns[3342] = 50'b10_0100100000111011_0100001001111100_0100000000111000;
      patterns[3343] = 50'b11_0100100000111011_0100001001111100_0100101001111111;
      patterns[3344] = 50'b00_0110010110101111_0110010101010110_1100101100000101;
      patterns[3345] = 50'b01_0110010110101111_0110010101010110_0000000001011001;
      patterns[3346] = 50'b10_0110010110101111_0110010101010110_0110010100000110;
      patterns[3347] = 50'b11_0110010110101111_0110010101010110_0110010111111111;
      patterns[3348] = 50'b00_0100001110111010_0100100011000010_1000110001111100;
      patterns[3349] = 50'b01_0100001110111010_0100100011000010_1111101011111000;
      patterns[3350] = 50'b10_0100001110111010_0100100011000010_0100000010000010;
      patterns[3351] = 50'b11_0100001110111010_0100100011000010_0100101111111010;
      patterns[3352] = 50'b00_1101010111001111_1110100001110010_1011111001000001;
      patterns[3353] = 50'b01_1101010111001111_1110100001110010_1110110101011101;
      patterns[3354] = 50'b10_1101010111001111_1110100001110010_1100000001000010;
      patterns[3355] = 50'b11_1101010111001111_1110100001110010_1111110111111111;
      patterns[3356] = 50'b00_0010100100100110_0011100111100011_0110001100001001;
      patterns[3357] = 50'b01_0010100100100110_0011100111100011_1110111101000011;
      patterns[3358] = 50'b10_0010100100100110_0011100111100011_0010100100100010;
      patterns[3359] = 50'b11_0010100100100110_0011100111100011_0011100111100111;
      patterns[3360] = 50'b00_0110011001011000_1100011100001011_0010110101100011;
      patterns[3361] = 50'b01_0110011001011000_1100011100001011_1001111101001101;
      patterns[3362] = 50'b10_0110011001011000_1100011100001011_0100011000001000;
      patterns[3363] = 50'b11_0110011001011000_1100011100001011_1110011101011011;
      patterns[3364] = 50'b00_1001101111110100_1000000000110001_0001110000100101;
      patterns[3365] = 50'b01_1001101111110100_1000000000110001_0001101111000011;
      patterns[3366] = 50'b10_1001101111110100_1000000000110001_1000000000110000;
      patterns[3367] = 50'b11_1001101111110100_1000000000110001_1001101111110101;
      patterns[3368] = 50'b00_1010001010011100_1001011010011111_0011100100111011;
      patterns[3369] = 50'b01_1010001010011100_1001011010011111_0000101111111101;
      patterns[3370] = 50'b10_1010001010011100_1001011010011111_1000001010011100;
      patterns[3371] = 50'b11_1010001010011100_1001011010011111_1011011010011111;
      patterns[3372] = 50'b00_0000001010010111_0101110001000001_0101111011011000;
      patterns[3373] = 50'b01_0000001010010111_0101110001000001_1010011001010110;
      patterns[3374] = 50'b10_0000001010010111_0101110001000001_0000000000000001;
      patterns[3375] = 50'b11_0000001010010111_0101110001000001_0101111011010111;
      patterns[3376] = 50'b00_1011001011010011_1101000100110000_1000010000000011;
      patterns[3377] = 50'b01_1011001011010011_1101000100110000_1110000110100011;
      patterns[3378] = 50'b10_1011001011010011_1101000100110000_1001000000010000;
      patterns[3379] = 50'b11_1011001011010011_1101000100110000_1111001111110011;
      patterns[3380] = 50'b00_1000001011011010_1110101001111011_0110110101010101;
      patterns[3381] = 50'b01_1000001011011010_1110101001111011_1001100001011111;
      patterns[3382] = 50'b10_1000001011011010_1110101001111011_1000001001011010;
      patterns[3383] = 50'b11_1000001011011010_1110101001111011_1110101011111011;
      patterns[3384] = 50'b00_1000100101111001_1101110100011010_0110011010010011;
      patterns[3385] = 50'b01_1000100101111001_1101110100011010_1010110001011111;
      patterns[3386] = 50'b10_1000100101111001_1101110100011010_1000100100011000;
      patterns[3387] = 50'b11_1000100101111001_1101110100011010_1101110101111011;
      patterns[3388] = 50'b00_1010001001010011_0010111110011110_1101000111110001;
      patterns[3389] = 50'b01_1010001001010011_0010111110011110_0111001010110101;
      patterns[3390] = 50'b10_1010001001010011_0010111110011110_0010001000010010;
      patterns[3391] = 50'b11_1010001001010011_0010111110011110_1010111111011111;
      patterns[3392] = 50'b00_1100101001001100_1101010000111100_1001111010001000;
      patterns[3393] = 50'b01_1100101001001100_1101010000111100_1111011000010000;
      patterns[3394] = 50'b10_1100101001001100_1101010000111100_1100000000001100;
      patterns[3395] = 50'b11_1100101001001100_1101010000111100_1101111001111100;
      patterns[3396] = 50'b00_1000011100100100_1001011011000100_0001110111101000;
      patterns[3397] = 50'b01_1000011100100100_1001011011000100_1111000001100000;
      patterns[3398] = 50'b10_1000011100100100_1001011011000100_1000011000000100;
      patterns[3399] = 50'b11_1000011100100100_1001011011000100_1001011111100100;
      patterns[3400] = 50'b00_1100111010000111_0011010110111100_0000010001000011;
      patterns[3401] = 50'b01_1100111010000111_0011010110111100_1001100011001011;
      patterns[3402] = 50'b10_1100111010000111_0011010110111100_0000010010000100;
      patterns[3403] = 50'b11_1100111010000111_0011010110111100_1111111110111111;
      patterns[3404] = 50'b00_0111111001011110_0011011011101000_1011010101000110;
      patterns[3405] = 50'b01_0111111001011110_0011011011101000_0100011101110110;
      patterns[3406] = 50'b10_0111111001011110_0011011011101000_0011011001001000;
      patterns[3407] = 50'b11_0111111001011110_0011011011101000_0111111011111110;
      patterns[3408] = 50'b00_0010011101101001_0000110011110011_0011010001011100;
      patterns[3409] = 50'b01_0010011101101001_0000110011110011_0001101001110110;
      patterns[3410] = 50'b10_0010011101101001_0000110011110011_0000010001100001;
      patterns[3411] = 50'b11_0010011101101001_0000110011110011_0010111111111011;
      patterns[3412] = 50'b00_1111111010010101_0100100100000111_0100011110011100;
      patterns[3413] = 50'b01_1111111010010101_0100100100000111_1011010110001110;
      patterns[3414] = 50'b10_1111111010010101_0100100100000111_0100100000000101;
      patterns[3415] = 50'b11_1111111010010101_0100100100000111_1111111110010111;
      patterns[3416] = 50'b00_0110010100111000_0001111101000100_1000010001111100;
      patterns[3417] = 50'b01_0110010100111000_0001111101000100_0100010111110100;
      patterns[3418] = 50'b10_0110010100111000_0001111101000100_0000010100000000;
      patterns[3419] = 50'b11_0110010100111000_0001111101000100_0111111101111100;
      patterns[3420] = 50'b00_1101011010010001_0111001101001110_0100100111011111;
      patterns[3421] = 50'b01_1101011010010001_0111001101001110_0110001101000011;
      patterns[3422] = 50'b10_1101011010010001_0111001101001110_0101001000000000;
      patterns[3423] = 50'b11_1101011010010001_0111001101001110_1111011111011111;
      patterns[3424] = 50'b00_1011011000111010_0110000111101001_0001100000100011;
      patterns[3425] = 50'b01_1011011000111010_0110000111101001_0101010001010001;
      patterns[3426] = 50'b10_1011011000111010_0110000111101001_0010000000101000;
      patterns[3427] = 50'b11_1011011000111010_0110000111101001_1111011111111011;
      patterns[3428] = 50'b00_1001100100100000_1111000100000011_1000101000100011;
      patterns[3429] = 50'b01_1001100100100000_1111000100000011_1010100000011101;
      patterns[3430] = 50'b10_1001100100100000_1111000100000011_1001000100000000;
      patterns[3431] = 50'b11_1001100100100000_1111000100000011_1111100100100011;
      patterns[3432] = 50'b00_0010011001100111_0101000000001110_0111011001110101;
      patterns[3433] = 50'b01_0010011001100111_0101000000001110_1101011001011001;
      patterns[3434] = 50'b10_0010011001100111_0101000000001110_0000000000000110;
      patterns[3435] = 50'b11_0010011001100111_0101000000001110_0111011001101111;
      patterns[3436] = 50'b00_1010000001111110_0010101000000110_1100101010000100;
      patterns[3437] = 50'b01_1010000001111110_0010101000000110_0111011001111000;
      patterns[3438] = 50'b10_1010000001111110_0010101000000110_0010000000000110;
      patterns[3439] = 50'b11_1010000001111110_0010101000000110_1010101001111110;
      patterns[3440] = 50'b00_1110010110111111_1011100010101011_1001111001101010;
      patterns[3441] = 50'b01_1110010110111111_1011100010101011_0010110100010100;
      patterns[3442] = 50'b10_1110010110111111_1011100010101011_1010000010101011;
      patterns[3443] = 50'b11_1110010110111111_1011100010101011_1111110110111111;
      patterns[3444] = 50'b00_0011010011010010_0000000000100011_0011010011110101;
      patterns[3445] = 50'b01_0011010011010010_0000000000100011_0011010010101111;
      patterns[3446] = 50'b10_0011010011010010_0000000000100011_0000000000000010;
      patterns[3447] = 50'b11_0011010011010010_0000000000100011_0011010011110011;
      patterns[3448] = 50'b00_0000000010001010_0100001100000001_0100001110001011;
      patterns[3449] = 50'b01_0000000010001010_0100001100000001_1011110110001001;
      patterns[3450] = 50'b10_0000000010001010_0100001100000001_0000000000000000;
      patterns[3451] = 50'b11_0000000010001010_0100001100000001_0100001110001011;
      patterns[3452] = 50'b00_0111101010101100_1111001110010010_0110111000111110;
      patterns[3453] = 50'b01_0111101010101100_1111001110010010_1000011100011010;
      patterns[3454] = 50'b10_0111101010101100_1111001110010010_0111001010000000;
      patterns[3455] = 50'b11_0111101010101100_1111001110010010_1111101110111110;
      patterns[3456] = 50'b00_0110000111111101_0011011110101011_1001100110101000;
      patterns[3457] = 50'b01_0110000111111101_0011011110101011_0010101001010010;
      patterns[3458] = 50'b10_0110000111111101_0011011110101011_0010000110101001;
      patterns[3459] = 50'b11_0110000111111101_0011011110101011_0111011111111111;
      patterns[3460] = 50'b00_1100111110011010_0100001101010111_0001001011110001;
      patterns[3461] = 50'b01_1100111110011010_0100001101010111_1000110001000011;
      patterns[3462] = 50'b10_1100111110011010_0100001101010111_0100001100010010;
      patterns[3463] = 50'b11_1100111110011010_0100001101010111_1100111111011111;
      patterns[3464] = 50'b00_1100111011101111_0001001110101001_1110001010011000;
      patterns[3465] = 50'b01_1100111011101111_0001001110101001_1011101101000110;
      patterns[3466] = 50'b10_1100111011101111_0001001110101001_0000001010101001;
      patterns[3467] = 50'b11_1100111011101111_0001001110101001_1101111111101111;
      patterns[3468] = 50'b00_0010010000100110_0101100101101101_0111110110010011;
      patterns[3469] = 50'b01_0010010000100110_0101100101101101_1100101010111001;
      patterns[3470] = 50'b10_0010010000100110_0101100101101101_0000000000100100;
      patterns[3471] = 50'b11_0010010000100110_0101100101101101_0111110101101111;
      patterns[3472] = 50'b00_1100001110101101_0000100111010010_1100110101111111;
      patterns[3473] = 50'b01_1100001110101101_0000100111010010_1011100111011011;
      patterns[3474] = 50'b10_1100001110101101_0000100111010010_0000000110000000;
      patterns[3475] = 50'b11_1100001110101101_0000100111010010_1100101111111111;
      patterns[3476] = 50'b00_1011001111100011_0010010111011110_1101100111000001;
      patterns[3477] = 50'b01_1011001111100011_0010010111011110_1000111000000101;
      patterns[3478] = 50'b10_1011001111100011_0010010111011110_0010000111000010;
      patterns[3479] = 50'b11_1011001111100011_0010010111011110_1011011111111111;
      patterns[3480] = 50'b00_1100010100010100_1101111010001101_1010001110100001;
      patterns[3481] = 50'b01_1100010100010100_1101111010001101_1110011010000111;
      patterns[3482] = 50'b10_1100010100010100_1101111010001101_1100010000000100;
      patterns[3483] = 50'b11_1100010100010100_1101111010001101_1101111110011101;
      patterns[3484] = 50'b00_0011010101011100_1000011100111001_1011110010010101;
      patterns[3485] = 50'b01_0011010101011100_1000011100111001_1010111000100011;
      patterns[3486] = 50'b10_0011010101011100_1000011100111001_0000010100011000;
      patterns[3487] = 50'b11_0011010101011100_1000011100111001_1011011101111101;
      patterns[3488] = 50'b00_1100001001111010_0111100011001111_0011101101001001;
      patterns[3489] = 50'b01_1100001001111010_0111100011001111_0100100110101011;
      patterns[3490] = 50'b10_1100001001111010_0111100011001111_0100000001001010;
      patterns[3491] = 50'b11_1100001001111010_0111100011001111_1111101011111111;
      patterns[3492] = 50'b00_0011110011111101_1000001000001101_1011111100001010;
      patterns[3493] = 50'b01_0011110011111101_1000001000001101_1011101011110000;
      patterns[3494] = 50'b10_0011110011111101_1000001000001101_0000000000001101;
      patterns[3495] = 50'b11_0011110011111101_1000001000001101_1011111011111101;
      patterns[3496] = 50'b00_1001101100010001_0001101010110001_1011010111000010;
      patterns[3497] = 50'b01_1001101100010001_0001101010110001_1000000001100000;
      patterns[3498] = 50'b10_1001101100010001_0001101010110001_0001101000010001;
      patterns[3499] = 50'b11_1001101100010001_0001101010110001_1001101110110001;
      patterns[3500] = 50'b00_0001011101011011_1101010001010110_1110101110110001;
      patterns[3501] = 50'b01_0001011101011011_1101010001010110_0100001100000101;
      patterns[3502] = 50'b10_0001011101011011_1101010001010110_0001010001010010;
      patterns[3503] = 50'b11_0001011101011011_1101010001010110_1101011101011111;
      patterns[3504] = 50'b00_1011011011010010_0111001100011001_0010100111101011;
      patterns[3505] = 50'b01_1011011011010010_0111001100011001_0100001110111001;
      patterns[3506] = 50'b10_1011011011010010_0111001100011001_0011001000010000;
      patterns[3507] = 50'b11_1011011011010010_0111001100011001_1111011111011011;
      patterns[3508] = 50'b00_1101000001100010_0110010100000001_0011010101100011;
      patterns[3509] = 50'b01_1101000001100010_0110010100000001_0110101101100001;
      patterns[3510] = 50'b10_1101000001100010_0110010100000001_0100000000000000;
      patterns[3511] = 50'b11_1101000001100010_0110010100000001_1111010101100011;
      patterns[3512] = 50'b00_1110100000010100_1010000101010100_1000100101101000;
      patterns[3513] = 50'b01_1110100000010100_1010000101010100_0100011011000000;
      patterns[3514] = 50'b10_1110100000010100_1010000101010100_1010000000010100;
      patterns[3515] = 50'b11_1110100000010100_1010000101010100_1110100101010100;
      patterns[3516] = 50'b00_0111011001011010_0010101011110011_1010000101001101;
      patterns[3517] = 50'b01_0111011001011010_0010101011110011_0100101101100111;
      patterns[3518] = 50'b10_0111011001011010_0010101011110011_0010001001010010;
      patterns[3519] = 50'b11_0111011001011010_0010101011110011_0111111011111011;
      patterns[3520] = 50'b00_0111100001010110_1101001010011110_0100101011110100;
      patterns[3521] = 50'b01_0111100001010110_1101001010011110_1010010110111000;
      patterns[3522] = 50'b10_0111100001010110_1101001010011110_0101000000010110;
      patterns[3523] = 50'b11_0111100001010110_1101001010011110_1111101011011110;
      patterns[3524] = 50'b00_1110100011001000_0110101001000110_0101001100001110;
      patterns[3525] = 50'b01_1110100011001000_0110101001000110_0111111010000010;
      patterns[3526] = 50'b10_1110100011001000_0110101001000110_0110100001000000;
      patterns[3527] = 50'b11_1110100011001000_0110101001000110_1110101011001110;
      patterns[3528] = 50'b00_0101011111110110_0101100011011110_1011000011010100;
      patterns[3529] = 50'b01_0101011111110110_0101100011011110_1111111100011000;
      patterns[3530] = 50'b10_0101011111110110_0101100011011110_0101000011010110;
      patterns[3531] = 50'b11_0101011111110110_0101100011011110_0101111111111110;
      patterns[3532] = 50'b00_1010110010010101_1001000110010000_0011111000100101;
      patterns[3533] = 50'b01_1010110010010101_1001000110010000_0001101100000101;
      patterns[3534] = 50'b10_1010110010010101_1001000110010000_1000000010010000;
      patterns[3535] = 50'b11_1010110010010101_1001000110010000_1011110110010101;
      patterns[3536] = 50'b00_1110010111001100_1111100100110001_1101111011111101;
      patterns[3537] = 50'b01_1110010111001100_1111100100110001_1110110010011011;
      patterns[3538] = 50'b10_1110010111001100_1111100100110001_1110000100000000;
      patterns[3539] = 50'b11_1110010111001100_1111100100110001_1111110111111101;
      patterns[3540] = 50'b00_0101000000001010_1001010001111001_1110010010000011;
      patterns[3541] = 50'b01_0101000000001010_1001010001111001_1011101110010001;
      patterns[3542] = 50'b10_0101000000001010_1001010001111001_0001000000001000;
      patterns[3543] = 50'b11_0101000000001010_1001010001111001_1101010001111011;
      patterns[3544] = 50'b00_1010100011011110_1011011111111111_0110000011011101;
      patterns[3545] = 50'b01_1010100011011110_1011011111111111_1111000011011111;
      patterns[3546] = 50'b10_1010100011011110_1011011111111111_1010000011011110;
      patterns[3547] = 50'b11_1010100011011110_1011011111111111_1011111111111111;
      patterns[3548] = 50'b00_1110001010000010_0101101111110101_0011111001110111;
      patterns[3549] = 50'b01_1110001010000010_0101101111110101_1000011010001101;
      patterns[3550] = 50'b10_1110001010000010_0101101111110101_0100001010000000;
      patterns[3551] = 50'b11_1110001010000010_0101101111110101_1111101111110111;
      patterns[3552] = 50'b00_1010001110110101_1001011110100101_0011101101011010;
      patterns[3553] = 50'b01_1010001110110101_1001011110100101_0000110000010000;
      patterns[3554] = 50'b10_1010001110110101_1001011110100101_1000001110100101;
      patterns[3555] = 50'b11_1010001110110101_1001011110100101_1011011110110101;
      patterns[3556] = 50'b00_1110010011100111_1100011111010111_1010110010111110;
      patterns[3557] = 50'b01_1110010011100111_1100011111010111_0001110100010000;
      patterns[3558] = 50'b10_1110010011100111_1100011111010111_1100010011000111;
      patterns[3559] = 50'b11_1110010011100111_1100011111010111_1110011111110111;
      patterns[3560] = 50'b00_1001110111111100_1001011000001010_0011010000000110;
      patterns[3561] = 50'b01_1001110111111100_1001011000001010_0000011111110010;
      patterns[3562] = 50'b10_1001110111111100_1001011000001010_1001010000001000;
      patterns[3563] = 50'b11_1001110111111100_1001011000001010_1001111111111110;
      patterns[3564] = 50'b00_1110000101010111_1100100010100001_1010100111111000;
      patterns[3565] = 50'b01_1110000101010111_1100100010100001_0001100010110110;
      patterns[3566] = 50'b10_1110000101010111_1100100010100001_1100000000000001;
      patterns[3567] = 50'b11_1110000101010111_1100100010100001_1110100111110111;
      patterns[3568] = 50'b00_1101111001110000_1011010010011010_1001001100001010;
      patterns[3569] = 50'b01_1101111001110000_1011010010011010_0010100111010110;
      patterns[3570] = 50'b10_1101111001110000_1011010010011010_1001010000010000;
      patterns[3571] = 50'b11_1101111001110000_1011010010011010_1111111011111010;
      patterns[3572] = 50'b00_1000100110001111_0100101111000010_1101010101010001;
      patterns[3573] = 50'b01_1000100110001111_0100101111000010_0011110111001101;
      patterns[3574] = 50'b10_1000100110001111_0100101111000010_0000100110000010;
      patterns[3575] = 50'b11_1000100110001111_0100101111000010_1100101111001111;
      patterns[3576] = 50'b00_0101010001010110_1111110101111100_0101000111010010;
      patterns[3577] = 50'b01_0101010001010110_1111110101111100_0101011011011010;
      patterns[3578] = 50'b10_0101010001010110_1111110101111100_0101010001010100;
      patterns[3579] = 50'b11_0101010001010110_1111110101111100_1111110101111110;
      patterns[3580] = 50'b00_1101010011100111_0000111110100101_1110010010001100;
      patterns[3581] = 50'b01_1101010011100111_0000111110100101_1100010101000010;
      patterns[3582] = 50'b10_1101010011100111_0000111110100101_0000010010100101;
      patterns[3583] = 50'b11_1101010011100111_0000111110100101_1101111111100111;
      patterns[3584] = 50'b00_0001110011110000_0100100000000101_0110010011110101;
      patterns[3585] = 50'b01_0001110011110000_0100100000000101_1101010011101011;
      patterns[3586] = 50'b10_0001110011110000_0100100000000101_0000100000000000;
      patterns[3587] = 50'b11_0001110011110000_0100100000000101_0101110011110101;
      patterns[3588] = 50'b00_0001100000001101_1111100000111101_0001000001001010;
      patterns[3589] = 50'b01_0001100000001101_1111100000111101_0001111111010000;
      patterns[3590] = 50'b10_0001100000001101_1111100000111101_0001100000001101;
      patterns[3591] = 50'b11_0001100000001101_1111100000111101_1111100000111101;
      patterns[3592] = 50'b00_1010011010101100_1111010110111011_1001110001100111;
      patterns[3593] = 50'b01_1010011010101100_1111010110111011_1011000011110001;
      patterns[3594] = 50'b10_1010011010101100_1111010110111011_1010010010101000;
      patterns[3595] = 50'b11_1010011010101100_1111010110111011_1111011110111111;
      patterns[3596] = 50'b00_0111100111001100_0010011111111010_1010000111000110;
      patterns[3597] = 50'b01_0111100111001100_0010011111111010_0101000111010010;
      patterns[3598] = 50'b10_0111100111001100_0010011111111010_0010000111001000;
      patterns[3599] = 50'b11_0111100111001100_0010011111111010_0111111111111110;
      patterns[3600] = 50'b00_0111000100001010_0000000001100111_0111000101110001;
      patterns[3601] = 50'b01_0111000100001010_0000000001100111_0111000010100011;
      patterns[3602] = 50'b10_0111000100001010_0000000001100111_0000000000000010;
      patterns[3603] = 50'b11_0111000100001010_0000000001100111_0111000101101111;
      patterns[3604] = 50'b00_0111100101111011_1111010001010011_0110110111001110;
      patterns[3605] = 50'b01_0111100101111011_1111010001010011_1000010100101000;
      patterns[3606] = 50'b10_0111100101111011_1111010001010011_0111000001010011;
      patterns[3607] = 50'b11_0111100101111011_1111010001010011_1111110101111011;
      patterns[3608] = 50'b00_1000110101101011_0111100100001001_0000011001110100;
      patterns[3609] = 50'b01_1000110101101011_0111100100001001_0001010001100010;
      patterns[3610] = 50'b10_1000110101101011_0111100100001001_0000100100001001;
      patterns[3611] = 50'b11_1000110101101011_0111100100001001_1111110101101011;
      patterns[3612] = 50'b00_0111010011110000_1100100001000110_0011110100110110;
      patterns[3613] = 50'b01_0111010011110000_1100100001000110_1010110010101010;
      patterns[3614] = 50'b10_0111010011110000_1100100001000110_0100000001000000;
      patterns[3615] = 50'b11_0111010011110000_1100100001000110_1111110011110110;
      patterns[3616] = 50'b00_1001001001010001_0000011010111000_1001100100001001;
      patterns[3617] = 50'b01_1001001001010001_0000011010111000_1000101110011001;
      patterns[3618] = 50'b10_1001001001010001_0000011010111000_0000001000010000;
      patterns[3619] = 50'b11_1001001001010001_0000011010111000_1001011011111001;
      patterns[3620] = 50'b00_0011110100010001_0010101010000000_0110011110010001;
      patterns[3621] = 50'b01_0011110100010001_0010101010000000_0001001010010001;
      patterns[3622] = 50'b10_0011110100010001_0010101010000000_0010100000000000;
      patterns[3623] = 50'b11_0011110100010001_0010101010000000_0011111110010001;
      patterns[3624] = 50'b00_1010011110111000_0000101110101011_1011001101100011;
      patterns[3625] = 50'b01_1010011110111000_0000101110101011_1001110000001101;
      patterns[3626] = 50'b10_1010011110111000_0000101110101011_0000001110101000;
      patterns[3627] = 50'b11_1010011110111000_0000101110101011_1010111110111011;
      patterns[3628] = 50'b00_1101000101011101_0110100000011001_0011100101110110;
      patterns[3629] = 50'b01_1101000101011101_0110100000011001_0110100101000100;
      patterns[3630] = 50'b10_1101000101011101_0110100000011001_0100000000011001;
      patterns[3631] = 50'b11_1101000101011101_0110100000011001_1111100101011101;
      patterns[3632] = 50'b00_1011000010010000_1101011000001010_1000011010011010;
      patterns[3633] = 50'b01_1011000010010000_1101011000001010_1101101010000110;
      patterns[3634] = 50'b10_1011000010010000_1101011000001010_1001000000000000;
      patterns[3635] = 50'b11_1011000010010000_1101011000001010_1111011010011010;
      patterns[3636] = 50'b00_0100110000000101_1101100000000010_0010010000000111;
      patterns[3637] = 50'b01_0100110000000101_1101100000000010_0111010000000011;
      patterns[3638] = 50'b10_0100110000000101_1101100000000010_0100100000000000;
      patterns[3639] = 50'b11_0100110000000101_1101100000000010_1101110000000111;
      patterns[3640] = 50'b00_0101101010001110_1010100101000000_0000001111001110;
      patterns[3641] = 50'b01_0101101010001110_1010100101000000_1011000101001110;
      patterns[3642] = 50'b10_0101101010001110_1010100101000000_0000100000000000;
      patterns[3643] = 50'b11_0101101010001110_1010100101000000_1111101111001110;
      patterns[3644] = 50'b00_1110000101110000_0100011010011101_0010100000001101;
      patterns[3645] = 50'b01_1110000101110000_0100011010011101_1001101011010011;
      patterns[3646] = 50'b10_1110000101110000_0100011010011101_0100000000010000;
      patterns[3647] = 50'b11_1110000101110000_0100011010011101_1110011111111101;
      patterns[3648] = 50'b00_0000101011001100_0111101111011100_1000011010101000;
      patterns[3649] = 50'b01_0000101011001100_0111101111011100_1000111011110000;
      patterns[3650] = 50'b10_0000101011001100_0111101111011100_0000101011001100;
      patterns[3651] = 50'b11_0000101011001100_0111101111011100_0111101111011100;
      patterns[3652] = 50'b00_1001011101000011_1101110000100010_0111001101100101;
      patterns[3653] = 50'b01_1001011101000011_1101110000100010_1011101100100001;
      patterns[3654] = 50'b10_1001011101000011_1101110000100010_1001010000000010;
      patterns[3655] = 50'b11_1001011101000011_1101110000100010_1101111101100011;
      patterns[3656] = 50'b00_0011001011110001_1111110101010010_0011000001000011;
      patterns[3657] = 50'b01_0011001011110001_1111110101010010_0011010110011111;
      patterns[3658] = 50'b10_0011001011110001_1111110101010010_0011000001010000;
      patterns[3659] = 50'b11_0011001011110001_1111110101010010_1111111111110011;
      patterns[3660] = 50'b00_0000000001001110_1011101110111000_1011110000000110;
      patterns[3661] = 50'b01_0000000001001110_1011101110111000_0100010010010110;
      patterns[3662] = 50'b10_0000000001001110_1011101110111000_0000000000001000;
      patterns[3663] = 50'b11_0000000001001110_1011101110111000_1011101111111110;
      patterns[3664] = 50'b00_1001011111100010_1101011000100000_0110111000000010;
      patterns[3665] = 50'b01_1001011111100010_1101011000100000_1100000111000010;
      patterns[3666] = 50'b10_1001011111100010_1101011000100000_1001011000100000;
      patterns[3667] = 50'b11_1001011111100010_1101011000100000_1101011111100010;
      patterns[3668] = 50'b00_1101101111101111_1010110001110100_1000100001100011;
      patterns[3669] = 50'b01_1101101111101111_1010110001110100_0010111101111011;
      patterns[3670] = 50'b10_1101101111101111_1010110001110100_1000100001100100;
      patterns[3671] = 50'b11_1101101111101111_1010110001110100_1111111111111111;
      patterns[3672] = 50'b00_0111100000110000_0001110000011011_1001010001001011;
      patterns[3673] = 50'b01_0111100000110000_0001110000011011_0101110000010101;
      patterns[3674] = 50'b10_0111100000110000_0001110000011011_0001100000010000;
      patterns[3675] = 50'b11_0111100000110000_0001110000011011_0111110000111011;
      patterns[3676] = 50'b00_1111000011000010_0101100010100011_0100100101100101;
      patterns[3677] = 50'b01_1111000011000010_0101100010100011_1001100000011111;
      patterns[3678] = 50'b10_1111000011000010_0101100010100011_0101000010000010;
      patterns[3679] = 50'b11_1111000011000010_0101100010100011_1111100011100011;
      patterns[3680] = 50'b00_0100110110111000_1010001111111101_1111000110110101;
      patterns[3681] = 50'b01_0100110110111000_1010001111111101_1010100110111011;
      patterns[3682] = 50'b10_0100110110111000_1010001111111101_0000000110111000;
      patterns[3683] = 50'b11_0100110110111000_1010001111111101_1110111111111101;
      patterns[3684] = 50'b00_1101101111001001_0001001100000110_1110111011001111;
      patterns[3685] = 50'b01_1101101111001001_0001001100000110_1100100011000011;
      patterns[3686] = 50'b10_1101101111001001_0001001100000110_0001001100000000;
      patterns[3687] = 50'b11_1101101111001001_0001001100000110_1101101111001111;
      patterns[3688] = 50'b00_0001101101000011_0011000001110100_0100101110110111;
      patterns[3689] = 50'b01_0001101101000011_0011000001110100_1110101011001111;
      patterns[3690] = 50'b10_0001101101000011_0011000001110100_0001000001000000;
      patterns[3691] = 50'b11_0001101101000011_0011000001110100_0011101101110111;
      patterns[3692] = 50'b00_1101011001011000_1001110011110101_0111001101001101;
      patterns[3693] = 50'b01_1101011001011000_1001110011110101_0011100101100011;
      patterns[3694] = 50'b10_1101011001011000_1001110011110101_1001010001010000;
      patterns[3695] = 50'b11_1101011001011000_1001110011110101_1101111011111101;
      patterns[3696] = 50'b00_1101010000000000_0111111000111001_0101001000111001;
      patterns[3697] = 50'b01_1101010000000000_0111111000111001_0101010111000111;
      patterns[3698] = 50'b10_1101010000000000_0111111000111001_0101010000000000;
      patterns[3699] = 50'b11_1101010000000000_0111111000111001_1111111000111001;
      patterns[3700] = 50'b00_1010011001011011_0001101110000101_1100000111100000;
      patterns[3701] = 50'b01_1010011001011011_0001101110000101_1000101011010110;
      patterns[3702] = 50'b10_1010011001011011_0001101110000101_0000001000000001;
      patterns[3703] = 50'b11_1010011001011011_0001101110000101_1011111111011111;
      patterns[3704] = 50'b00_0111000000110111_1101010000000101_0100010000111100;
      patterns[3705] = 50'b01_0111000000110111_1101010000000101_1001110000110010;
      patterns[3706] = 50'b10_0111000000110111_1101010000000101_0101000000000101;
      patterns[3707] = 50'b11_0111000000110111_1101010000000101_1111010000110111;
      patterns[3708] = 50'b00_0000010111100010_0100010100100101_0100101100000111;
      patterns[3709] = 50'b01_0000010111100010_0100010100100101_1100000010111101;
      patterns[3710] = 50'b10_0000010111100010_0100010100100101_0000010100100000;
      patterns[3711] = 50'b11_0000010111100010_0100010100100101_0100010111100111;
      patterns[3712] = 50'b00_1010111110001101_0000110001100010_1011101111101111;
      patterns[3713] = 50'b01_1010111110001101_0000110001100010_1010001100101011;
      patterns[3714] = 50'b10_1010111110001101_0000110001100010_0000110000000000;
      patterns[3715] = 50'b11_1010111110001101_0000110001100010_1010111111101111;
      patterns[3716] = 50'b00_1100111111111011_1101010001011001_1010010001010100;
      patterns[3717] = 50'b01_1100111111111011_1101010001011001_1111101110100010;
      patterns[3718] = 50'b10_1100111111111011_1101010001011001_1100010001011001;
      patterns[3719] = 50'b11_1100111111111011_1101010001011001_1101111111111011;
      patterns[3720] = 50'b00_0101111010101111_0000011010100100_0110010101010011;
      patterns[3721] = 50'b01_0101111010101111_0000011010100100_0101100000001011;
      patterns[3722] = 50'b10_0101111010101111_0000011010100100_0000011010100100;
      patterns[3723] = 50'b11_0101111010101111_0000011010100100_0101111010101111;
      patterns[3724] = 50'b00_0010101001000000_0111011101111010_1010000110111010;
      patterns[3725] = 50'b01_0010101001000000_0111011101111010_1011001011000110;
      patterns[3726] = 50'b10_0010101001000000_0111011101111010_0010001001000000;
      patterns[3727] = 50'b11_0010101001000000_0111011101111010_0111111101111010;
      patterns[3728] = 50'b00_0011001101000101_0000101110100010_0011111011100111;
      patterns[3729] = 50'b01_0011001101000101_0000101110100010_0010011110100011;
      patterns[3730] = 50'b10_0011001101000101_0000101110100010_0000001100000000;
      patterns[3731] = 50'b11_0011001101000101_0000101110100010_0011101111100111;
      patterns[3732] = 50'b00_1011001110101001_1100100010101111_0111110001011000;
      patterns[3733] = 50'b01_1011001110101001_1100100010101111_1110101011111010;
      patterns[3734] = 50'b10_1011001110101001_1100100010101111_1000000010101001;
      patterns[3735] = 50'b11_1011001110101001_1100100010101111_1111101110101111;
      patterns[3736] = 50'b00_1111011001111100_1111100111100010_1111000001011110;
      patterns[3737] = 50'b01_1111011001111100_1111100111100010_1111110010011010;
      patterns[3738] = 50'b10_1111011001111100_1111100111100010_1111000001100000;
      patterns[3739] = 50'b11_1111011001111100_1111100111100010_1111111111111110;
      patterns[3740] = 50'b00_0111101010000111_0101010001110110_1100111011111101;
      patterns[3741] = 50'b01_0111101010000111_0101010001110110_0010011000010001;
      patterns[3742] = 50'b10_0111101010000111_0101010001110110_0101000000000110;
      patterns[3743] = 50'b11_0111101010000111_0101010001110110_0111111011110111;
      patterns[3744] = 50'b00_1100001110011001_1111110001010001_1011111111101010;
      patterns[3745] = 50'b01_1100001110011001_1111110001010001_1100011101001000;
      patterns[3746] = 50'b10_1100001110011001_1111110001010001_1100000000010001;
      patterns[3747] = 50'b11_1100001110011001_1111110001010001_1111111111011001;
      patterns[3748] = 50'b00_0001110010111000_0101100001111111_0111010100110111;
      patterns[3749] = 50'b01_0001110010111000_0101100001111111_1100010000111001;
      patterns[3750] = 50'b10_0001110010111000_0101100001111111_0001100000111000;
      patterns[3751] = 50'b11_0001110010111000_0101100001111111_0101110011111111;
      patterns[3752] = 50'b00_1001010101000110_0010010111010101_1011101100011011;
      patterns[3753] = 50'b01_1001010101000110_0010010111010101_0110111101110001;
      patterns[3754] = 50'b10_1001010101000110_0010010111010101_0000010101000100;
      patterns[3755] = 50'b11_1001010101000110_0010010111010101_1011010111010111;
      patterns[3756] = 50'b00_1111111001110101_1010111110101110_1010111000100011;
      patterns[3757] = 50'b01_1111111001110101_1010111110101110_0100111011000111;
      patterns[3758] = 50'b10_1111111001110101_1010111110101110_1010111000100100;
      patterns[3759] = 50'b11_1111111001110101_1010111110101110_1111111111111111;
      patterns[3760] = 50'b00_0011100110100010_1000101100110000_1100010011010010;
      patterns[3761] = 50'b01_0011100110100010_1000101100110000_1010111001110010;
      patterns[3762] = 50'b10_0011100110100010_1000101100110000_0000100100100000;
      patterns[3763] = 50'b11_0011100110100010_1000101100110000_1011101110110010;
      patterns[3764] = 50'b00_1111010101010000_0101001101111011_0100100011001011;
      patterns[3765] = 50'b01_1111010101010000_0101001101111011_1010000111010101;
      patterns[3766] = 50'b10_1111010101010000_0101001101111011_0101000101010000;
      patterns[3767] = 50'b11_1111010101010000_0101001101111011_1111011101111011;
      patterns[3768] = 50'b00_0000101001000111_0101110000010011_0110011001011010;
      patterns[3769] = 50'b01_0000101001000111_0101110000010011_1010111000110100;
      patterns[3770] = 50'b10_0000101001000111_0101110000010011_0000100000000011;
      patterns[3771] = 50'b11_0000101001000111_0101110000010011_0101111001010111;
      patterns[3772] = 50'b00_0001111000111101_1111011000011000_0001010001010101;
      patterns[3773] = 50'b01_0001111000111101_1111011000011000_0010100000100101;
      patterns[3774] = 50'b10_0001111000111101_1111011000011000_0001011000011000;
      patterns[3775] = 50'b11_0001111000111101_1111011000011000_1111111000111101;
      patterns[3776] = 50'b00_0111001010111110_0000101101100000_0111111000011110;
      patterns[3777] = 50'b01_0111001010111110_0000101101100000_0110011101011110;
      patterns[3778] = 50'b10_0111001010111110_0000101101100000_0000001000100000;
      patterns[3779] = 50'b11_0111001010111110_0000101101100000_0111101111111110;
      patterns[3780] = 50'b00_1101011011000011_0111101111111101_0101001011000000;
      patterns[3781] = 50'b01_1101011011000011_0111101111111101_0101101011000110;
      patterns[3782] = 50'b10_1101011011000011_0111101111111101_0101001011000001;
      patterns[3783] = 50'b11_1101011011000011_0111101111111101_1111111111111111;
      patterns[3784] = 50'b00_0110010100100000_1100110111011111_0011001011111111;
      patterns[3785] = 50'b01_0110010100100000_1100110111011111_1001011101000001;
      patterns[3786] = 50'b10_0110010100100000_1100110111011111_0100010100000000;
      patterns[3787] = 50'b11_0110010100100000_1100110111011111_1110110111111111;
      patterns[3788] = 50'b00_1111101010100110_1000011011010100_1000000101111010;
      patterns[3789] = 50'b01_1111101010100110_1000011011010100_0111001111010010;
      patterns[3790] = 50'b10_1111101010100110_1000011011010100_1000001010000100;
      patterns[3791] = 50'b11_1111101010100110_1000011011010100_1111111011110110;
      patterns[3792] = 50'b00_0101100111010111_1001011000001001_1110111111100000;
      patterns[3793] = 50'b01_0101100111010111_1001011000001001_1100001111001110;
      patterns[3794] = 50'b10_0101100111010111_1001011000001001_0001000000000001;
      patterns[3795] = 50'b11_0101100111010111_1001011000001001_1101111111011111;
      patterns[3796] = 50'b00_1001100010110110_1101011011100011_0110111110011001;
      patterns[3797] = 50'b01_1001100010110110_1101011011100011_1100000111010011;
      patterns[3798] = 50'b10_1001100010110110_1101011011100011_1001000010100010;
      patterns[3799] = 50'b11_1001100010110110_1101011011100011_1101111011110111;
      patterns[3800] = 50'b00_0101110011000000_0011101010001011_1001011101001011;
      patterns[3801] = 50'b01_0101110011000000_0011101010001011_0010001000110101;
      patterns[3802] = 50'b10_0101110011000000_0011101010001011_0001100010000000;
      patterns[3803] = 50'b11_0101110011000000_0011101010001011_0111111011001011;
      patterns[3804] = 50'b00_0100101001111111_0000001101011111_0100110111011110;
      patterns[3805] = 50'b01_0100101001111111_0000001101011111_0100011100100000;
      patterns[3806] = 50'b10_0100101001111111_0000001101011111_0000001001011111;
      patterns[3807] = 50'b11_0100101001111111_0000001101011111_0100101101111111;
      patterns[3808] = 50'b00_1111011100101001_1010010010111000_1001101111100001;
      patterns[3809] = 50'b01_1111011100101001_1010010010111000_0101001001110001;
      patterns[3810] = 50'b10_1111011100101001_1010010010111000_1010010000101000;
      patterns[3811] = 50'b11_1111011100101001_1010010010111000_1111011110111001;
      patterns[3812] = 50'b00_0011110000011101_1110110101011111_0010100101111100;
      patterns[3813] = 50'b01_0011110000011101_1110110101011111_0100111010111110;
      patterns[3814] = 50'b10_0011110000011101_1110110101011111_0010110000011101;
      patterns[3815] = 50'b11_0011110000011101_1110110101011111_1111110101011111;
      patterns[3816] = 50'b00_0111101101011001_1011101100001101_0011011001100110;
      patterns[3817] = 50'b01_0111101101011001_1011101100001101_1100000001001100;
      patterns[3818] = 50'b10_0111101101011001_1011101100001101_0011101100001001;
      patterns[3819] = 50'b11_0111101101011001_1011101100001101_1111101101011101;
      patterns[3820] = 50'b00_1011101001100010_0101110001000000_0001011010100010;
      patterns[3821] = 50'b01_1011101001100010_0101110001000000_0101111000100010;
      patterns[3822] = 50'b10_1011101001100010_0101110001000000_0001100001000000;
      patterns[3823] = 50'b11_1011101001100010_0101110001000000_1111111001100010;
      patterns[3824] = 50'b00_0101001110101101_0011101101101110_1000111100011011;
      patterns[3825] = 50'b01_0101001110101101_0011101101101110_0001100000111111;
      patterns[3826] = 50'b10_0101001110101101_0011101101101110_0001001100101100;
      patterns[3827] = 50'b11_0101001110101101_0011101101101110_0111101111101111;
      patterns[3828] = 50'b00_1100111100001100_0110010111000000_0011010011001100;
      patterns[3829] = 50'b01_1100111100001100_0110010111000000_0110100101001100;
      patterns[3830] = 50'b10_1100111100001100_0110010111000000_0100010100000000;
      patterns[3831] = 50'b11_1100111100001100_0110010111000000_1110111111001100;
      patterns[3832] = 50'b00_0111110001110011_1101111111001110_0101110001000001;
      patterns[3833] = 50'b01_0111110001110011_1101111111001110_1001110010100101;
      patterns[3834] = 50'b10_0111110001110011_1101111111001110_0101110001000010;
      patterns[3835] = 50'b11_0111110001110011_1101111111001110_1111111111111111;
      patterns[3836] = 50'b00_0000101111010001_1001111100100110_1010101011110111;
      patterns[3837] = 50'b01_0000101111010001_1001111100100110_0110110010101011;
      patterns[3838] = 50'b10_0000101111010001_1001111100100110_0000101100000000;
      patterns[3839] = 50'b11_0000101111010001_1001111100100110_1001111111110111;
      patterns[3840] = 50'b00_0011110100001101_1111011101100101_0011010001110010;
      patterns[3841] = 50'b01_0011110100001101_1111011101100101_0100010110101000;
      patterns[3842] = 50'b10_0011110100001101_1111011101100101_0011010100000101;
      patterns[3843] = 50'b11_0011110100001101_1111011101100101_1111111101101101;
      patterns[3844] = 50'b00_0010011001011110_1001100000100111_1011111010000101;
      patterns[3845] = 50'b01_0010011001011110_1001100000100111_1000111000110111;
      patterns[3846] = 50'b10_0010011001011110_1001100000100111_0000000000000110;
      patterns[3847] = 50'b11_0010011001011110_1001100000100111_1011111001111111;
      patterns[3848] = 50'b00_1000101000001010_0001010110100011_1001111110101101;
      patterns[3849] = 50'b01_1000101000001010_0001010110100011_0111010001100111;
      patterns[3850] = 50'b10_1000101000001010_0001010110100011_0000000000000010;
      patterns[3851] = 50'b11_1000101000001010_0001010110100011_1001111110101011;
      patterns[3852] = 50'b00_0111000010101000_1100101101111011_0011110000100011;
      patterns[3853] = 50'b01_0111000010101000_1100101101111011_1010010100101101;
      patterns[3854] = 50'b10_0111000010101000_1100101101111011_0100000000101000;
      patterns[3855] = 50'b11_0111000010101000_1100101101111011_1111101111111011;
      patterns[3856] = 50'b00_0011011100110010_1001011110000111_1100111010111001;
      patterns[3857] = 50'b01_0011011100110010_1001011110000111_1001111110101011;
      patterns[3858] = 50'b10_0011011100110010_1001011110000111_0001011100000010;
      patterns[3859] = 50'b11_0011011100110010_1001011110000111_1011011110110111;
      patterns[3860] = 50'b00_1000101000101010_0000010000110111_1000111001100001;
      patterns[3861] = 50'b01_1000101000101010_0000010000110111_1000010111110011;
      patterns[3862] = 50'b10_1000101000101010_0000010000110111_0000000000100010;
      patterns[3863] = 50'b11_1000101000101010_0000010000110111_1000111000111111;
      patterns[3864] = 50'b00_0100010111000101_1000011100000011_1100110011001000;
      patterns[3865] = 50'b01_0100010111000101_1000011100000011_1011111011000010;
      patterns[3866] = 50'b10_0100010111000101_1000011100000011_0000010100000001;
      patterns[3867] = 50'b11_0100010111000101_1000011100000011_1100011111000111;
      patterns[3868] = 50'b00_1101111111011011_0011001001101110_0001001001001001;
      patterns[3869] = 50'b01_1101111111011011_0011001001101110_1010110101101101;
      patterns[3870] = 50'b10_1101111111011011_0011001001101110_0001001001001010;
      patterns[3871] = 50'b11_1101111111011011_0011001001101110_1111111111111111;
      patterns[3872] = 50'b00_0010100001100000_1101001110011100_1111101111111100;
      patterns[3873] = 50'b01_0010100001100000_1101001110011100_0101010011000100;
      patterns[3874] = 50'b10_0010100001100000_1101001110011100_0000000000000000;
      patterns[3875] = 50'b11_0010100001100000_1101001110011100_1111101111111100;
      patterns[3876] = 50'b00_1011001000010001_1100110010110100_0111111011000101;
      patterns[3877] = 50'b01_1011001000010001_1100110010110100_1110010101011101;
      patterns[3878] = 50'b10_1011001000010001_1100110010110100_1000000000010000;
      patterns[3879] = 50'b11_1011001000010001_1100110010110100_1111111010110101;
      patterns[3880] = 50'b00_1100101101000010_1110111001101011_1011100110101101;
      patterns[3881] = 50'b01_1100101101000010_1110111001101011_1101110011010111;
      patterns[3882] = 50'b10_1100101101000010_1110111001101011_1100101001000010;
      patterns[3883] = 50'b11_1100101101000010_1110111001101011_1110111101101011;
      patterns[3884] = 50'b00_0110000010001110_0010011101101101_1000011111111011;
      patterns[3885] = 50'b01_0110000010001110_0010011101101101_0011100100100001;
      patterns[3886] = 50'b10_0110000010001110_0010011101101101_0010000000001100;
      patterns[3887] = 50'b11_0110000010001110_0010011101101101_0110011111101111;
      patterns[3888] = 50'b00_1000110011101111_1001011100101010_0010010000011001;
      patterns[3889] = 50'b01_1000110011101111_1001011100101010_1111010111000101;
      patterns[3890] = 50'b10_1000110011101111_1001011100101010_1000010000101010;
      patterns[3891] = 50'b11_1000110011101111_1001011100101010_1001111111101111;
      patterns[3892] = 50'b00_1010111001100010_1001111000011100_0100110001111110;
      patterns[3893] = 50'b01_1010111001100010_1001111000011100_0001000001000110;
      patterns[3894] = 50'b10_1010111001100010_1001111000011100_1000111000000000;
      patterns[3895] = 50'b11_1010111001100010_1001111000011100_1011111001111110;
      patterns[3896] = 50'b00_0001100001101111_0000111011111010_0010011101101001;
      patterns[3897] = 50'b01_0001100001101111_0000111011111010_0000100101110101;
      patterns[3898] = 50'b10_0001100001101111_0000111011111010_0000100001101010;
      patterns[3899] = 50'b11_0001100001101111_0000111011111010_0001111011111111;
      patterns[3900] = 50'b00_1000100010000000_0000011000010010_1000111010010010;
      patterns[3901] = 50'b01_1000100010000000_0000011000010010_1000001001101110;
      patterns[3902] = 50'b10_1000100010000000_0000011000010010_0000000000000000;
      patterns[3903] = 50'b11_1000100010000000_0000011000010010_1000111010010010;
      patterns[3904] = 50'b00_0011111110010000_1111010100001000_0011010010011000;
      patterns[3905] = 50'b01_0011111110010000_1111010100001000_0100101010001000;
      patterns[3906] = 50'b10_0011111110010000_1111010100001000_0011010100000000;
      patterns[3907] = 50'b11_0011111110010000_1111010100001000_1111111110011000;
      patterns[3908] = 50'b00_1001101100001011_1010010100101100_0100000000110111;
      patterns[3909] = 50'b01_1001101100001011_1010010100101100_1111010111011111;
      patterns[3910] = 50'b10_1001101100001011_1010010100101100_1000000100001000;
      patterns[3911] = 50'b11_1001101100001011_1010010100101100_1011111100101111;
      patterns[3912] = 50'b00_1000100100000001_1100100000111110_0101000100111111;
      patterns[3913] = 50'b01_1000100100000001_1100100000111110_1100000011000011;
      patterns[3914] = 50'b10_1000100100000001_1100100000111110_1000100000000000;
      patterns[3915] = 50'b11_1000100100000001_1100100000111110_1100100100111111;
      patterns[3916] = 50'b00_1010101011001110_1101001010001001_0111110101010111;
      patterns[3917] = 50'b01_1010101011001110_1101001010001001_1101100001000101;
      patterns[3918] = 50'b10_1010101011001110_1101001010001001_1000001010001000;
      patterns[3919] = 50'b11_1010101011001110_1101001010001001_1111101011001111;
      patterns[3920] = 50'b00_0010001100100111_0110100010100111_1000101111001110;
      patterns[3921] = 50'b01_0010001100100111_0110100010100111_1011101010000000;
      patterns[3922] = 50'b10_0010001100100111_0110100010100111_0010000000100111;
      patterns[3923] = 50'b11_0010001100100111_0110100010100111_0110101110100111;
      patterns[3924] = 50'b00_0011100101100100_0111101001100001_1011001111000101;
      patterns[3925] = 50'b01_0011100101100100_0111101001100001_1011111100000011;
      patterns[3926] = 50'b10_0011100101100100_0111101001100001_0011100001100000;
      patterns[3927] = 50'b11_0011100101100100_0111101001100001_0111101101100101;
      patterns[3928] = 50'b00_0101000111110110_1111101000110111_0100110000101101;
      patterns[3929] = 50'b01_0101000111110110_1111101000110111_0101011110111111;
      patterns[3930] = 50'b10_0101000111110110_1111101000110111_0101000000110110;
      patterns[3931] = 50'b11_0101000111110110_1111101000110111_1111101111110111;
      patterns[3932] = 50'b00_0111001111111101_1111100101101000_0110110101100101;
      patterns[3933] = 50'b01_0111001111111101_1111100101101000_0111101010010101;
      patterns[3934] = 50'b10_0111001111111101_1111100101101000_0111000101101000;
      patterns[3935] = 50'b11_0111001111111101_1111100101101000_1111101111111101;
      patterns[3936] = 50'b00_0011101100111111_0011101000010000_0111010101001111;
      patterns[3937] = 50'b01_0011101100111111_0011101000010000_0000000100101111;
      patterns[3938] = 50'b10_0011101100111111_0011101000010000_0011101000010000;
      patterns[3939] = 50'b11_0011101100111111_0011101000010000_0011101100111111;
      patterns[3940] = 50'b00_1100110111001000_0010011101100111_1111010100101111;
      patterns[3941] = 50'b01_1100110111001000_0010011101100111_1010011001100001;
      patterns[3942] = 50'b10_1100110111001000_0010011101100111_0000010101000000;
      patterns[3943] = 50'b11_1100110111001000_0010011101100111_1110111111101111;
      patterns[3944] = 50'b00_0010101000110010_1010111010001101_1101100010111111;
      patterns[3945] = 50'b01_0010101000110010_1010111010001101_0111101110100101;
      patterns[3946] = 50'b10_0010101000110010_1010111010001101_0010101000000000;
      patterns[3947] = 50'b11_0010101000110010_1010111010001101_1010111010111111;
      patterns[3948] = 50'b00_1111000001101001_1111001111110111_1110010001100000;
      patterns[3949] = 50'b01_1111000001101001_1111001111110111_1111110001110010;
      patterns[3950] = 50'b10_1111000001101001_1111001111110111_1111000001100001;
      patterns[3951] = 50'b11_1111000001101001_1111001111110111_1111001111111111;
      patterns[3952] = 50'b00_0000000000001011_0001100110010010_0001100110011101;
      patterns[3953] = 50'b01_0000000000001011_0001100110010010_1110011001111001;
      patterns[3954] = 50'b10_0000000000001011_0001100110010010_0000000000000010;
      patterns[3955] = 50'b11_0000000000001011_0001100110010010_0001100110011011;
      patterns[3956] = 50'b00_1101111000001101_1010101110000000_1000100110001101;
      patterns[3957] = 50'b01_1101111000001101_1010101110000000_0011001010001101;
      patterns[3958] = 50'b10_1101111000001101_1010101110000000_1000101000000000;
      patterns[3959] = 50'b11_1101111000001101_1010101110000000_1111111110001101;
      patterns[3960] = 50'b00_1000110100101001_0011101111111011_1100100100100100;
      patterns[3961] = 50'b01_1000110100101001_0011101111111011_0101000100101110;
      patterns[3962] = 50'b10_1000110100101001_0011101111111011_0000100100101001;
      patterns[3963] = 50'b11_1000110100101001_0011101111111011_1011111111111011;
      patterns[3964] = 50'b00_0011100111111101_1101010111110010_0000111111101111;
      patterns[3965] = 50'b01_0011100111111101_1101010111110010_0110010000001011;
      patterns[3966] = 50'b10_0011100111111101_1101010111110010_0001000111110000;
      patterns[3967] = 50'b11_0011100111111101_1101010111110010_1111110111111111;
      patterns[3968] = 50'b00_1111101011111111_0100100000100111_0100001100100110;
      patterns[3969] = 50'b01_1111101011111111_0100100000100111_1011001011011000;
      patterns[3970] = 50'b10_1111101011111111_0100100000100111_0100100000100111;
      patterns[3971] = 50'b11_1111101011111111_0100100000100111_1111101011111111;
      patterns[3972] = 50'b00_1010110111000011_1010001111011010_0101000110011101;
      patterns[3973] = 50'b01_1010110111000011_1010001111011010_0000100111101001;
      patterns[3974] = 50'b10_1010110111000011_1010001111011010_1010000111000010;
      patterns[3975] = 50'b11_1010110111000011_1010001111011010_1010111111011011;
      patterns[3976] = 50'b00_0100010010100100_0101100011101101_1001110110010001;
      patterns[3977] = 50'b01_0100010010100100_0101100011101101_1110101110110111;
      patterns[3978] = 50'b10_0100010010100100_0101100011101101_0100000010100100;
      patterns[3979] = 50'b11_0100010010100100_0101100011101101_0101110011101101;
      patterns[3980] = 50'b00_0100101000111111_0000100110111011_0101001111111010;
      patterns[3981] = 50'b01_0100101000111111_0000100110111011_0100000010000100;
      patterns[3982] = 50'b10_0100101000111111_0000100110111011_0000100000111011;
      patterns[3983] = 50'b11_0100101000111111_0000100110111011_0100101110111111;
      patterns[3984] = 50'b00_1111100011111010_1110000110001100_1101101010000110;
      patterns[3985] = 50'b01_1111100011111010_1110000110001100_0001011101101110;
      patterns[3986] = 50'b10_1111100011111010_1110000110001100_1110000010001000;
      patterns[3987] = 50'b11_1111100011111010_1110000110001100_1111100111111110;
      patterns[3988] = 50'b00_1001010101001100_1111110011100001_1001001000101101;
      patterns[3989] = 50'b01_1001010101001100_1111110011100001_1001100001101011;
      patterns[3990] = 50'b10_1001010101001100_1111110011100001_1001010001000000;
      patterns[3991] = 50'b11_1001010101001100_1111110011100001_1111110111101101;
      patterns[3992] = 50'b00_0010011010010111_0101001001010001_0111100011101000;
      patterns[3993] = 50'b01_0010011010010111_0101001001010001_1101010001000110;
      patterns[3994] = 50'b10_0010011010010111_0101001001010001_0000001000010001;
      patterns[3995] = 50'b11_0010011010010111_0101001001010001_0111011011010111;
      patterns[3996] = 50'b00_1010110110111000_1100000000000100_0110110110111100;
      patterns[3997] = 50'b01_1010110110111000_1100000000000100_1110110110110100;
      patterns[3998] = 50'b10_1010110110111000_1100000000000100_1000000000000000;
      patterns[3999] = 50'b11_1010110110111000_1100000000000100_1110110110111100;
      patterns[4000] = 50'b00_0101111100001001_0001110100001110_0111110000010111;
      patterns[4001] = 50'b01_0101111100001001_0001110100001110_0100000111111011;
      patterns[4002] = 50'b10_0101111100001001_0001110100001110_0001110100001000;
      patterns[4003] = 50'b11_0101111100001001_0001110100001110_0101111100001111;
      patterns[4004] = 50'b00_1001000011001110_1101000101111101_0110001001001011;
      patterns[4005] = 50'b01_1001000011001110_1101000101111101_1011111101010001;
      patterns[4006] = 50'b10_1001000011001110_1101000101111101_1001000001001100;
      patterns[4007] = 50'b11_1001000011001110_1101000101111101_1101000111111111;
      patterns[4008] = 50'b00_0011010000001000_1101101110011111_0000111110100111;
      patterns[4009] = 50'b01_0011010000001000_1101101110011111_0101100001101001;
      patterns[4010] = 50'b10_0011010000001000_1101101110011111_0001000000001000;
      patterns[4011] = 50'b11_0011010000001000_1101101110011111_1111111110011111;
      patterns[4012] = 50'b00_0001010110100111_1101011111100100_1110110110001011;
      patterns[4013] = 50'b01_0001010110100111_1101011111100100_0011110111000011;
      patterns[4014] = 50'b10_0001010110100111_1101011111100100_0001010110100100;
      patterns[4015] = 50'b11_0001010110100111_1101011111100100_1101011111100111;
      patterns[4016] = 50'b00_0110111010110111_1001101000001100_0000100011000011;
      patterns[4017] = 50'b01_0110111010110111_1001101000001100_1101010010101011;
      patterns[4018] = 50'b10_0110111010110111_1001101000001100_0000101000000100;
      patterns[4019] = 50'b11_0110111010110111_1001101000001100_1111111010111111;
      patterns[4020] = 50'b00_1010001111110010_1101110101001001_1000000100111011;
      patterns[4021] = 50'b01_1010001111110010_1101110101001001_1100011010101001;
      patterns[4022] = 50'b10_1010001111110010_1101110101001001_1000000101000000;
      patterns[4023] = 50'b11_1010001111110010_1101110101001001_1111111111111011;
      patterns[4024] = 50'b00_1000011000001110_0010110100010100_1011001100100010;
      patterns[4025] = 50'b01_1000011000001110_0010110100010100_0101100011111010;
      patterns[4026] = 50'b10_1000011000001110_0010110100010100_0000010000000100;
      patterns[4027] = 50'b11_1000011000001110_0010110100010100_1010111100011110;
      patterns[4028] = 50'b00_0000010100001100_0100010001101111_0100100101111011;
      patterns[4029] = 50'b01_0000010100001100_0100010001101111_1100000010011101;
      patterns[4030] = 50'b10_0000010100001100_0100010001101111_0000010000001100;
      patterns[4031] = 50'b11_0000010100001100_0100010001101111_0100010101101111;
      patterns[4032] = 50'b00_1000011011111001_0000110100100111_1001010000100000;
      patterns[4033] = 50'b01_1000011011111001_0000110100100111_0111100111010010;
      patterns[4034] = 50'b10_1000011011111001_0000110100100111_0000010000100001;
      patterns[4035] = 50'b11_1000011011111001_0000110100100111_1000111111111111;
      patterns[4036] = 50'b00_1110111101110100_0010011010111011_0001011000101111;
      patterns[4037] = 50'b01_1110111101110100_0010011010111011_1100100010111001;
      patterns[4038] = 50'b10_1110111101110100_0010011010111011_0010011000110000;
      patterns[4039] = 50'b11_1110111101110100_0010011010111011_1110111111111111;
      patterns[4040] = 50'b00_1011010111100100_0110010100011100_0001101100000000;
      patterns[4041] = 50'b01_1011010111100100_0110010100011100_0101000011001000;
      patterns[4042] = 50'b10_1011010111100100_0110010100011100_0010010100000100;
      patterns[4043] = 50'b11_1011010111100100_0110010100011100_1111010111111100;
      patterns[4044] = 50'b00_0001011000001000_0011010010110010_0100101010111010;
      patterns[4045] = 50'b01_0001011000001000_0011010010110010_1110000101010110;
      patterns[4046] = 50'b10_0001011000001000_0011010010110010_0001010000000000;
      patterns[4047] = 50'b11_0001011000001000_0011010010110010_0011011010111010;
      patterns[4048] = 50'b00_1010111010100101_1110001100101101_1001000111010010;
      patterns[4049] = 50'b01_1010111010100101_1110001100101101_1100101101111000;
      patterns[4050] = 50'b10_1010111010100101_1110001100101101_1010001000100101;
      patterns[4051] = 50'b11_1010111010100101_1110001100101101_1110111110101101;
      patterns[4052] = 50'b00_1001010110010011_1100011001000001_0101101111010100;
      patterns[4053] = 50'b01_1001010110010011_1100011001000001_1100111101010010;
      patterns[4054] = 50'b10_1001010110010011_1100011001000001_1000010000000001;
      patterns[4055] = 50'b11_1001010110010011_1100011001000001_1101011111010011;
      patterns[4056] = 50'b00_1010110100001101_0110000111111011_0000111100001000;
      patterns[4057] = 50'b01_1010110100001101_0110000111111011_0100101100010010;
      patterns[4058] = 50'b10_1010110100001101_0110000111111011_0010000100001001;
      patterns[4059] = 50'b11_1010110100001101_0110000111111011_1110110111111111;
      patterns[4060] = 50'b00_1001010010010010_1000001100101101_0001011110111111;
      patterns[4061] = 50'b01_1001010010010010_1000001100101101_0001000101100101;
      patterns[4062] = 50'b10_1001010010010010_1000001100101101_1000000000000000;
      patterns[4063] = 50'b11_1001010010010010_1000001100101101_1001011110111111;
      patterns[4064] = 50'b00_1111010110000111_1010111010110110_1010010000111101;
      patterns[4065] = 50'b01_1111010110000111_1010111010110110_0100011011010001;
      patterns[4066] = 50'b10_1111010110000111_1010111010110110_1010010010000110;
      patterns[4067] = 50'b11_1111010110000111_1010111010110110_1111111110110111;
      patterns[4068] = 50'b00_1100101001001001_1110111101010110_1011100110011111;
      patterns[4069] = 50'b01_1100101001001001_1110111101010110_1101101011110011;
      patterns[4070] = 50'b10_1100101001001001_1110111101010110_1100101001000000;
      patterns[4071] = 50'b11_1100101001001001_1110111101010110_1110111101011111;
      patterns[4072] = 50'b00_0000101010010010_1000100010011110_1001001100110000;
      patterns[4073] = 50'b01_0000101010010010_1000100010011110_1000000111110100;
      patterns[4074] = 50'b10_0000101010010010_1000100010011110_0000100010010010;
      patterns[4075] = 50'b11_0000101010010010_1000100010011110_1000101010011110;
      patterns[4076] = 50'b00_0110101101111001_0011000110111111_1001110100111000;
      patterns[4077] = 50'b01_0110101101111001_0011000110111111_0011100110111010;
      patterns[4078] = 50'b10_0110101101111001_0011000110111111_0010000100111001;
      patterns[4079] = 50'b11_0110101101111001_0011000110111111_0111101111111111;
      patterns[4080] = 50'b00_0111100100000001_0111010101110100_1110111001110101;
      patterns[4081] = 50'b01_0111100100000001_0111010101110100_0000001110001101;
      patterns[4082] = 50'b10_0111100100000001_0111010101110100_0111000100000000;
      patterns[4083] = 50'b11_0111100100000001_0111010101110100_0111110101110101;
      patterns[4084] = 50'b00_1010110001011101_1010000010000001_0100110011011110;
      patterns[4085] = 50'b01_1010110001011101_1010000010000001_0000101111011100;
      patterns[4086] = 50'b10_1010110001011101_1010000010000001_1010000000000001;
      patterns[4087] = 50'b11_1010110001011101_1010000010000001_1010110011011101;
      patterns[4088] = 50'b00_1000101001001000_0010110110100101_1011011111101101;
      patterns[4089] = 50'b01_1000101001001000_0010110110100101_0101110010100011;
      patterns[4090] = 50'b10_1000101001001000_0010110110100101_0000100000000000;
      patterns[4091] = 50'b11_1000101001001000_0010110110100101_1010111111101101;
      patterns[4092] = 50'b00_1010000011000001_1111011100000111_1001011111001000;
      patterns[4093] = 50'b01_1010000011000001_1111011100000111_1010100110111010;
      patterns[4094] = 50'b10_1010000011000001_1111011100000111_1010000000000001;
      patterns[4095] = 50'b11_1010000011000001_1111011100000111_1111011111000111;
      patterns[4096] = 50'b00_0001100101000010_0011001000110100_0100101101110110;
      patterns[4097] = 50'b01_0001100101000010_0011001000110100_1110011100001110;
      patterns[4098] = 50'b10_0001100101000010_0011001000110100_0001000000000000;
      patterns[4099] = 50'b11_0001100101000010_0011001000110100_0011101101110110;
      patterns[4100] = 50'b00_1100010001001010_1001111101010101_0110001110011111;
      patterns[4101] = 50'b01_1100010001001010_1001111101010101_0010010011110101;
      patterns[4102] = 50'b10_1100010001001010_1001111101010101_1000010001000000;
      patterns[4103] = 50'b11_1100010001001010_1001111101010101_1101111101011111;
      patterns[4104] = 50'b00_0001101100111001_1001010110101000_1011000011100001;
      patterns[4105] = 50'b01_0001101100111001_1001010110101000_1000010110010001;
      patterns[4106] = 50'b10_0001101100111001_1001010110101000_0001000100101000;
      patterns[4107] = 50'b11_0001101100111001_1001010110101000_1001111110111001;
      patterns[4108] = 50'b00_1101111001010100_0010001000110000_0000000010000100;
      patterns[4109] = 50'b01_1101111001010100_0010001000110000_1011110000100100;
      patterns[4110] = 50'b10_1101111001010100_0010001000110000_0000001000010000;
      patterns[4111] = 50'b11_1101111001010100_0010001000110000_1111111001110100;
      patterns[4112] = 50'b00_0010110000011000_0010000010011011_0100110010110011;
      patterns[4113] = 50'b01_0010110000011000_0010000010011011_0000101101111101;
      patterns[4114] = 50'b10_0010110000011000_0010000010011011_0010000000011000;
      patterns[4115] = 50'b11_0010110000011000_0010000010011011_0010110010011011;
      patterns[4116] = 50'b00_0100010111110100_1010010101011000_1110101101001100;
      patterns[4117] = 50'b01_0100010111110100_1010010101011000_1010000010011100;
      patterns[4118] = 50'b10_0100010111110100_1010010101011000_0000010101010000;
      patterns[4119] = 50'b11_0100010111110100_1010010101011000_1110010111111100;
      patterns[4120] = 50'b00_1001001000011000_1100000110100000_0101001110111000;
      patterns[4121] = 50'b01_1001001000011000_1100000110100000_1101000001111000;
      patterns[4122] = 50'b10_1001001000011000_1100000110100000_1000000000000000;
      patterns[4123] = 50'b11_1001001000011000_1100000110100000_1101001110111000;
      patterns[4124] = 50'b00_1100010000000000_0101101001000001_0001111001000001;
      patterns[4125] = 50'b01_1100010000000000_0101101001000001_0110100110111111;
      patterns[4126] = 50'b10_1100010000000000_0101101001000001_0100000000000000;
      patterns[4127] = 50'b11_1100010000000000_0101101001000001_1101111001000001;
      patterns[4128] = 50'b00_1011101001001001_1010011110010000_0110000111011001;
      patterns[4129] = 50'b01_1011101001001001_1010011110010000_0001001010111001;
      patterns[4130] = 50'b10_1011101001001001_1010011110010000_1010001000000000;
      patterns[4131] = 50'b11_1011101001001001_1010011110010000_1011111111011001;
      patterns[4132] = 50'b00_0111001000110110_1110001011101100_0101010100100010;
      patterns[4133] = 50'b01_0111001000110110_1110001011101100_1000111101001010;
      patterns[4134] = 50'b10_0111001000110110_1110001011101100_0110001000100100;
      patterns[4135] = 50'b11_0111001000110110_1110001011101100_1111001011111110;
      patterns[4136] = 50'b00_0010010011001000_0111110010010100_1010000101011100;
      patterns[4137] = 50'b01_0010010011001000_0111110010010100_1010100000110100;
      patterns[4138] = 50'b10_0010010011001000_0111110010010100_0010010010000000;
      patterns[4139] = 50'b11_0010010011001000_0111110010010100_0111110011011100;
      patterns[4140] = 50'b00_1111111111010100_1111110111010101_1111110110101001;
      patterns[4141] = 50'b01_1111111111010100_1111110111010101_0000000111111111;
      patterns[4142] = 50'b10_1111111111010100_1111110111010101_1111110111010100;
      patterns[4143] = 50'b11_1111111111010100_1111110111010101_1111111111010101;
      patterns[4144] = 50'b00_0001010010001010_1111011101011101_0000101111100111;
      patterns[4145] = 50'b01_0001010010001010_1111011101011101_0001110100101101;
      patterns[4146] = 50'b10_0001010010001010_1111011101011101_0001010000001000;
      patterns[4147] = 50'b11_0001010010001010_1111011101011101_1111011111011111;
      patterns[4148] = 50'b00_1011010101000111_0011110100011011_1111001001100010;
      patterns[4149] = 50'b01_1011010101000111_0011110100011011_0111100000101100;
      patterns[4150] = 50'b10_1011010101000111_0011110100011011_0011010100000011;
      patterns[4151] = 50'b11_1011010101000111_0011110100011011_1011110101011111;
      patterns[4152] = 50'b00_0001101111111110_0101111101110010_0111101101110000;
      patterns[4153] = 50'b01_0001101111111110_0101111101110010_1011110010001100;
      patterns[4154] = 50'b10_0001101111111110_0101111101110010_0001101101110010;
      patterns[4155] = 50'b11_0001101111111110_0101111101110010_0101111111111110;
      patterns[4156] = 50'b00_0110100111000101_0010100001000111_1001001000001100;
      patterns[4157] = 50'b01_0110100111000101_0010100001000111_0100000101111110;
      patterns[4158] = 50'b10_0110100111000101_0010100001000111_0010100001000101;
      patterns[4159] = 50'b11_0110100111000101_0010100001000111_0110100111000111;
      patterns[4160] = 50'b00_1100110100000101_1011000010000010_0111110110000111;
      patterns[4161] = 50'b01_1100110100000101_1011000010000010_0001110010000011;
      patterns[4162] = 50'b10_1100110100000101_1011000010000010_1000000000000000;
      patterns[4163] = 50'b11_1100110100000101_1011000010000010_1111110110000111;
      patterns[4164] = 50'b00_0101111011101000_1110101101101000_0100101001010000;
      patterns[4165] = 50'b01_0101111011101000_1110101101101000_0111001110000000;
      patterns[4166] = 50'b10_0101111011101000_1110101101101000_0100101001101000;
      patterns[4167] = 50'b11_0101111011101000_1110101101101000_1111111111101000;
      patterns[4168] = 50'b00_0110011111101110_1100000000011011_0010100000001001;
      patterns[4169] = 50'b01_0110011111101110_1100000000011011_1010011111010011;
      patterns[4170] = 50'b10_0110011111101110_1100000000011011_0100000000001010;
      patterns[4171] = 50'b11_0110011111101110_1100000000011011_1110011111111111;
      patterns[4172] = 50'b00_1001111110101111_1010000101011100_0100000100001011;
      patterns[4173] = 50'b01_1001111110101111_1010000101011100_1111111001010011;
      patterns[4174] = 50'b10_1001111110101111_1010000101011100_1000000100001100;
      patterns[4175] = 50'b11_1001111110101111_1010000101011100_1011111111111111;
      patterns[4176] = 50'b00_0110001001111000_0010100000111110_1000101010110110;
      patterns[4177] = 50'b01_0110001001111000_0010100000111110_0011101000111010;
      patterns[4178] = 50'b10_0110001001111000_0010100000111110_0010000000111000;
      patterns[4179] = 50'b11_0110001001111000_0010100000111110_0110101001111110;
      patterns[4180] = 50'b00_0001000101110001_0101101010001000_0110101111111001;
      patterns[4181] = 50'b01_0001000101110001_0101101010001000_1011011011101001;
      patterns[4182] = 50'b10_0001000101110001_0101101010001000_0001000000000000;
      patterns[4183] = 50'b11_0001000101110001_0101101010001000_0101101111111001;
      patterns[4184] = 50'b00_0000010100010101_1100000010100111_1100010110111100;
      patterns[4185] = 50'b01_0000010100010101_1100000010100111_0100010001101110;
      patterns[4186] = 50'b10_0000010100010101_1100000010100111_0000000000000101;
      patterns[4187] = 50'b11_0000010100010101_1100000010100111_1100010110110111;
      patterns[4188] = 50'b00_1101111010101010_0011110001010011_0001101011111101;
      patterns[4189] = 50'b01_1101111010101010_0011110001010011_1010001001010111;
      patterns[4190] = 50'b10_1101111010101010_0011110001010011_0001110000000010;
      patterns[4191] = 50'b11_1101111010101010_0011110001010011_1111111011111011;
      patterns[4192] = 50'b00_0010100111100010_0001111111001100_0100100110101110;
      patterns[4193] = 50'b01_0010100111100010_0001111111001100_0000101000010110;
      patterns[4194] = 50'b10_0010100111100010_0001111111001100_0000100111000000;
      patterns[4195] = 50'b11_0010100111100010_0001111111001100_0011111111101110;
      patterns[4196] = 50'b00_0100010010101111_0111100100010110_1011110111000101;
      patterns[4197] = 50'b01_0100010010101111_0111100100010110_1100101110011001;
      patterns[4198] = 50'b10_0100010010101111_0111100100010110_0100000000000110;
      patterns[4199] = 50'b11_0100010010101111_0111100100010110_0111110110111111;
      patterns[4200] = 50'b00_0101111000010011_1111001111011101_0101000111110000;
      patterns[4201] = 50'b01_0101111000010011_1111001111011101_0110101000110110;
      patterns[4202] = 50'b10_0101111000010011_1111001111011101_0101001000010001;
      patterns[4203] = 50'b11_0101111000010011_1111001111011101_1111111111011111;
      patterns[4204] = 50'b00_0001011010101110_0110101101110101_1000001000100011;
      patterns[4205] = 50'b01_0001011010101110_0110101101110101_1010101100111001;
      patterns[4206] = 50'b10_0001011010101110_0110101101110101_0000001000100100;
      patterns[4207] = 50'b11_0001011010101110_0110101101110101_0111111111111111;
      patterns[4208] = 50'b00_0100001111001001_0000001101010100_0100011100011101;
      patterns[4209] = 50'b01_0100001111001001_0000001101010100_0100000001110101;
      patterns[4210] = 50'b10_0100001111001001_0000001101010100_0000001101000000;
      patterns[4211] = 50'b11_0100001111001001_0000001101010100_0100001111011101;
      patterns[4212] = 50'b00_0111100110001111_1101001100110110_0100110011000101;
      patterns[4213] = 50'b01_0111100110001111_1101001100110110_1010011001011001;
      patterns[4214] = 50'b10_0111100110001111_1101001100110110_0101000100000110;
      patterns[4215] = 50'b11_0111100110001111_1101001100110110_1111101110111111;
      patterns[4216] = 50'b00_0001011110010100_0100101111011001_0110001101101101;
      patterns[4217] = 50'b01_0001011110010100_0100101111011001_1100101110111011;
      patterns[4218] = 50'b10_0001011110010100_0100101111011001_0000001110010000;
      patterns[4219] = 50'b11_0001011110010100_0100101111011001_0101111111011101;
      patterns[4220] = 50'b00_0111010110001110_0000110100010101_1000001010100011;
      patterns[4221] = 50'b01_0111010110001110_0000110100010101_0110100001111001;
      patterns[4222] = 50'b10_0111010110001110_0000110100010101_0000010100000100;
      patterns[4223] = 50'b11_0111010110001110_0000110100010101_0111110110011111;
      patterns[4224] = 50'b00_1010101000001110_0000010110001100_1010111110011010;
      patterns[4225] = 50'b01_1010101000001110_0000010110001100_1010010010000010;
      patterns[4226] = 50'b10_1010101000001110_0000010110001100_0000000000001100;
      patterns[4227] = 50'b11_1010101000001110_0000010110001100_1010111110001110;
      patterns[4228] = 50'b00_1111101110101010_0010001000110001_0001110111011011;
      patterns[4229] = 50'b01_1111101110101010_0010001000110001_1101100101111001;
      patterns[4230] = 50'b10_1111101110101010_0010001000110001_0010001000100000;
      patterns[4231] = 50'b11_1111101110101010_0010001000110001_1111101110111011;
      patterns[4232] = 50'b00_1111001101010111_0100011111101111_0011101101000110;
      patterns[4233] = 50'b01_1111001101010111_0100011111101111_1010101101101000;
      patterns[4234] = 50'b10_1111001101010111_0100011111101111_0100001101000111;
      patterns[4235] = 50'b11_1111001101010111_0100011111101111_1111011111111111;
      patterns[4236] = 50'b00_1110011001001000_1011011100000000_1001110101001000;
      patterns[4237] = 50'b01_1110011001001000_1011011100000000_0010111101001000;
      patterns[4238] = 50'b10_1110011001001000_1011011100000000_1010011000000000;
      patterns[4239] = 50'b11_1110011001001000_1011011100000000_1111011101001000;
      patterns[4240] = 50'b00_1010001101011110_1010110100010100_0101000001110010;
      patterns[4241] = 50'b01_1010001101011110_1010110100010100_1111011001001010;
      patterns[4242] = 50'b10_1010001101011110_1010110100010100_1010000100010100;
      patterns[4243] = 50'b11_1010001101011110_1010110100010100_1010111101011110;
      patterns[4244] = 50'b00_0100110110011001_0011010011111101_1000001010010110;
      patterns[4245] = 50'b01_0100110110011001_0011010011111101_0001100010011100;
      patterns[4246] = 50'b10_0100110110011001_0011010011111101_0000010010011001;
      patterns[4247] = 50'b11_0100110110011001_0011010011111101_0111110111111101;
      patterns[4248] = 50'b00_1011011101000000_1001011010111010_0100110111111010;
      patterns[4249] = 50'b01_1011011101000000_1001011010111010_0010000010000110;
      patterns[4250] = 50'b10_1011011101000000_1001011010111010_1001011000000000;
      patterns[4251] = 50'b11_1011011101000000_1001011010111010_1011011111111010;
      patterns[4252] = 50'b00_0100000110101000_0000010101100101_0100011100001101;
      patterns[4253] = 50'b01_0100000110101000_0000010101100101_0011110001000011;
      patterns[4254] = 50'b10_0100000110101000_0000010101100101_0000000100100000;
      patterns[4255] = 50'b11_0100000110101000_0000010101100101_0100010111101101;
      patterns[4256] = 50'b00_0010100100101100_1010100010000000_1101000110101100;
      patterns[4257] = 50'b01_0010100100101100_1010100010000000_1000000010101100;
      patterns[4258] = 50'b10_0010100100101100_1010100010000000_0010100000000000;
      patterns[4259] = 50'b11_0010100100101100_1010100010000000_1010100110101100;
      patterns[4260] = 50'b00_1001110100100011_0101011011000110_1111001111101001;
      patterns[4261] = 50'b01_1001110100100011_0101011011000110_0100011001011101;
      patterns[4262] = 50'b10_1001110100100011_0101011011000110_0001010000000010;
      patterns[4263] = 50'b11_1001110100100011_0101011011000110_1101111111100111;
      patterns[4264] = 50'b00_0100010110000110_1010000101100011_1110011011101001;
      patterns[4265] = 50'b01_0100010110000110_1010000101100011_1010010000100011;
      patterns[4266] = 50'b10_0100010110000110_1010000101100011_0000000100000010;
      patterns[4267] = 50'b11_0100010110000110_1010000101100011_1110010111100111;
      patterns[4268] = 50'b00_0010110100111101_1011001000110100_1101111101110001;
      patterns[4269] = 50'b01_0010110100111101_1011001000110100_0111101100001001;
      patterns[4270] = 50'b10_0010110100111101_1011001000110100_0010000000110100;
      patterns[4271] = 50'b11_0010110100111101_1011001000110100_1011111100111101;
      patterns[4272] = 50'b00_0000110101001100_1111111000011010_0000101101100110;
      patterns[4273] = 50'b01_0000110101001100_1111111000011010_0000111100110010;
      patterns[4274] = 50'b10_0000110101001100_1111111000011010_0000110000001000;
      patterns[4275] = 50'b11_0000110101001100_1111111000011010_1111111101011110;
      patterns[4276] = 50'b00_1101110000111111_1001100001011110_0111010010011101;
      patterns[4277] = 50'b01_1101110000111111_1001100001011110_0100001111100001;
      patterns[4278] = 50'b10_1101110000111111_1001100001011110_1001100000011110;
      patterns[4279] = 50'b11_1101110000111111_1001100001011110_1101110001111111;
      patterns[4280] = 50'b00_0101001011101101_1011010100011100_0000100000001001;
      patterns[4281] = 50'b01_0101001011101101_1011010100011100_1001110111010001;
      patterns[4282] = 50'b10_0101001011101101_1011010100011100_0001000000001100;
      patterns[4283] = 50'b11_0101001011101101_1011010100011100_1111011111111101;
      patterns[4284] = 50'b00_1110010110100110_0111100111100110_0101111110001100;
      patterns[4285] = 50'b01_1110010110100110_0111100111100110_0110101111000000;
      patterns[4286] = 50'b10_1110010110100110_0111100111100110_0110000110100110;
      patterns[4287] = 50'b11_1110010110100110_0111100111100110_1111110111100110;
      patterns[4288] = 50'b00_1110110000010011_1110110001010100_1101100001100111;
      patterns[4289] = 50'b01_1110110000010011_1110110001010100_1111111110111111;
      patterns[4290] = 50'b10_1110110000010011_1110110001010100_1110110000010000;
      patterns[4291] = 50'b11_1110110000010011_1110110001010100_1110110001010111;
      patterns[4292] = 50'b00_0101101111100110_1010000110100110_1111110110001100;
      patterns[4293] = 50'b01_0101101111100110_1010000110100110_1011101001000000;
      patterns[4294] = 50'b10_0101101111100110_1010000110100110_0000000110100110;
      patterns[4295] = 50'b11_0101101111100110_1010000110100110_1111101111100110;
      patterns[4296] = 50'b00_0110100000011000_1011111111001111_0010011111100111;
      patterns[4297] = 50'b01_0110100000011000_1011111111001111_1010100001001001;
      patterns[4298] = 50'b10_0110100000011000_1011111111001111_0010100000001000;
      patterns[4299] = 50'b11_0110100000011000_1011111111001111_1111111111011111;
      patterns[4300] = 50'b00_0111000100101110_0001001011001001_1000001111110111;
      patterns[4301] = 50'b01_0111000100101110_0001001011001001_0101111001100101;
      patterns[4302] = 50'b10_0111000100101110_0001001011001001_0001000000001000;
      patterns[4303] = 50'b11_0111000100101110_0001001011001001_0111001111101111;
      patterns[4304] = 50'b00_0011100000011001_0000111111110011_0100100000001100;
      patterns[4305] = 50'b01_0011100000011001_0000111111110011_0010100000100110;
      patterns[4306] = 50'b10_0011100000011001_0000111111110011_0000100000010001;
      patterns[4307] = 50'b11_0011100000011001_0000111111110011_0011111111111011;
      patterns[4308] = 50'b00_0000010111000000_1110111111101111_1111010110101111;
      patterns[4309] = 50'b01_0000010111000000_1110111111101111_0001010111010001;
      patterns[4310] = 50'b10_0000010111000000_1110111111101111_0000010111000000;
      patterns[4311] = 50'b11_0000010111000000_1110111111101111_1110111111101111;
      patterns[4312] = 50'b00_0001101011110001_1101010011111111_1110111111110000;
      patterns[4313] = 50'b01_0001101011110001_1101010011111111_0100010111110010;
      patterns[4314] = 50'b10_0001101011110001_1101010011111111_0001000011110001;
      patterns[4315] = 50'b11_0001101011110001_1101010011111111_1101111011111111;
      patterns[4316] = 50'b00_1111011111000011_1011101110110010_1011001101110101;
      patterns[4317] = 50'b01_1111011111000011_1011101110110010_0011110000010001;
      patterns[4318] = 50'b10_1111011111000011_1011101110110010_1011001110000010;
      patterns[4319] = 50'b11_1111011111000011_1011101110110010_1111111111110011;
      patterns[4320] = 50'b00_1110110010000101_1010010011101010_1001000101101111;
      patterns[4321] = 50'b01_1110110010000101_1010010011101010_0100011110011011;
      patterns[4322] = 50'b10_1110110010000101_1010010011101010_1010010010000000;
      patterns[4323] = 50'b11_1110110010000101_1010010011101010_1110110011101111;
      patterns[4324] = 50'b00_1001000110011110_1010011001001001_0011011111100111;
      patterns[4325] = 50'b01_1001000110011110_1010011001001001_1110101101010101;
      patterns[4326] = 50'b10_1001000110011110_1010011001001001_1000000000001000;
      patterns[4327] = 50'b11_1001000110011110_1010011001001001_1011011111011111;
      patterns[4328] = 50'b00_1010110100100100_1110111111011110_1001110100000010;
      patterns[4329] = 50'b01_1010110100100100_1110111111011110_1011110101000110;
      patterns[4330] = 50'b10_1010110100100100_1110111111011110_1010110100000100;
      patterns[4331] = 50'b11_1010110100100100_1110111111011110_1110111111111110;
      patterns[4332] = 50'b00_0011110100111001_0010011100100111_0110010001100000;
      patterns[4333] = 50'b01_0011110100111001_0010011100100111_0001011000010010;
      patterns[4334] = 50'b10_0011110100111001_0010011100100111_0010010100100001;
      patterns[4335] = 50'b11_0011110100111001_0010011100100111_0011111100111111;
      patterns[4336] = 50'b00_1011001011110100_1111011011101001_1010100111011101;
      patterns[4337] = 50'b01_1011001011110100_1111011011101001_1011110000001011;
      patterns[4338] = 50'b10_1011001011110100_1111011011101001_1011001011100000;
      patterns[4339] = 50'b11_1011001011110100_1111011011101001_1111011011111101;
      patterns[4340] = 50'b00_0101001111001001_0101010011000110_1010100010001111;
      patterns[4341] = 50'b01_0101001111001001_0101010011000110_1111111100000011;
      patterns[4342] = 50'b10_0101001111001001_0101010011000110_0101000011000000;
      patterns[4343] = 50'b11_0101001111001001_0101010011000110_0101011111001111;
      patterns[4344] = 50'b00_0111110010100110_1010011110011001_0010010000111111;
      patterns[4345] = 50'b01_0111110010100110_1010011110011001_1101010100001101;
      patterns[4346] = 50'b10_0111110010100110_1010011110011001_0010010010000000;
      patterns[4347] = 50'b11_0111110010100110_1010011110011001_1111111110111111;
      patterns[4348] = 50'b00_0111101011100111_1100100000000100_0100001011101011;
      patterns[4349] = 50'b01_0111101011100111_1100100000000100_1011001011100011;
      patterns[4350] = 50'b10_0111101011100111_1100100000000100_0100100000000100;
      patterns[4351] = 50'b11_0111101011100111_1100100000000100_1111101011100111;
      patterns[4352] = 50'b00_1000100111101100_0101011010100100_1110000010010000;
      patterns[4353] = 50'b01_1000100111101100_0101011010100100_0011001101001000;
      patterns[4354] = 50'b10_1000100111101100_0101011010100100_0000000010100100;
      patterns[4355] = 50'b11_1000100111101100_0101011010100100_1101111111101100;
      patterns[4356] = 50'b00_1000000100101011_0101101110111010_1101110011100101;
      patterns[4357] = 50'b01_1000000100101011_0101101110111010_0010010101110001;
      patterns[4358] = 50'b10_1000000100101011_0101101110111010_0000000100101010;
      patterns[4359] = 50'b11_1000000100101011_0101101110111010_1101101110111011;
      patterns[4360] = 50'b00_1111001101100000_1100101011010011_1011111000110011;
      patterns[4361] = 50'b01_1111001101100000_1100101011010011_0010100010001101;
      patterns[4362] = 50'b10_1111001101100000_1100101011010011_1100001001000000;
      patterns[4363] = 50'b11_1111001101100000_1100101011010011_1111101111110011;
      patterns[4364] = 50'b00_0001010110010010_1100010010001000_1101101000011010;
      patterns[4365] = 50'b01_0001010110010010_1100010010001000_0101000100001010;
      patterns[4366] = 50'b10_0001010110010010_1100010010001000_0000010010000000;
      patterns[4367] = 50'b11_0001010110010010_1100010010001000_1101010110011010;
      patterns[4368] = 50'b00_0011100011101110_0010100011001001_0110000110110111;
      patterns[4369] = 50'b01_0011100011101110_0010100011001001_0001000000100101;
      patterns[4370] = 50'b10_0011100011101110_0010100011001001_0010100011001000;
      patterns[4371] = 50'b11_0011100011101110_0010100011001001_0011100011101111;
      patterns[4372] = 50'b00_0000011001000111_1100111111100010_1101011000101001;
      patterns[4373] = 50'b01_0000011001000111_1100111111100010_0011011001100101;
      patterns[4374] = 50'b10_0000011001000111_1100111111100010_0000011001000010;
      patterns[4375] = 50'b11_0000011001000111_1100111111100010_1100111111100111;
      patterns[4376] = 50'b00_1110001011011110_0001011101011110_1111101000111100;
      patterns[4377] = 50'b01_1110001011011110_0001011101011110_1100101110000000;
      patterns[4378] = 50'b10_1110001011011110_0001011101011110_0000001001011110;
      patterns[4379] = 50'b11_1110001011011110_0001011101011110_1111011111011110;
      patterns[4380] = 50'b00_1110110010111000_0001010011100011_0000000110011011;
      patterns[4381] = 50'b01_1110110010111000_0001010011100011_1101011111010101;
      patterns[4382] = 50'b10_1110110010111000_0001010011100011_0000010010100000;
      patterns[4383] = 50'b11_1110110010111000_0001010011100011_1111110011111011;
      patterns[4384] = 50'b00_0001111100010001_1110001110101110_0000001010111111;
      patterns[4385] = 50'b01_0001111100010001_1110001110101110_0011101101100011;
      patterns[4386] = 50'b10_0001111100010001_1110001110101110_0000001100000000;
      patterns[4387] = 50'b11_0001111100010001_1110001110101110_1111111110111111;
      patterns[4388] = 50'b00_0100111000000011_0000010010000110_0101001010001001;
      patterns[4389] = 50'b01_0100111000000011_0000010010000110_0100100101111101;
      patterns[4390] = 50'b10_0100111000000011_0000010010000110_0000010000000010;
      patterns[4391] = 50'b11_0100111000000011_0000010010000110_0100111010000111;
      patterns[4392] = 50'b00_0111100100011010_1000001100011000_1111110000110010;
      patterns[4393] = 50'b01_0111100100011010_1000001100011000_1111011000000010;
      patterns[4394] = 50'b10_0111100100011010_1000001100011000_0000000100011000;
      patterns[4395] = 50'b11_0111100100011010_1000001100011000_1111101100011010;
      patterns[4396] = 50'b00_0100000000011101_1001001000101001_1101001001000110;
      patterns[4397] = 50'b01_0100000000011101_1001001000101001_1010110111110100;
      patterns[4398] = 50'b10_0100000000011101_1001001000101001_0000000000001001;
      patterns[4399] = 50'b11_0100000000011101_1001001000101001_1101001000111101;
      patterns[4400] = 50'b00_0010100100110111_0001000010110001_0011100111101000;
      patterns[4401] = 50'b01_0010100100110111_0001000010110001_0001100010000110;
      patterns[4402] = 50'b10_0010100100110111_0001000010110001_0000000000110001;
      patterns[4403] = 50'b11_0010100100110111_0001000010110001_0011100110110111;
      patterns[4404] = 50'b00_1001010101001001_0010000010010010_1011010111011011;
      patterns[4405] = 50'b01_1001010101001001_0010000010010010_0111010010110111;
      patterns[4406] = 50'b10_1001010101001001_0010000010010010_0000000000000000;
      patterns[4407] = 50'b11_1001010101001001_0010000010010010_1011010111011011;
      patterns[4408] = 50'b00_0011101101011101_1100101100001101_0000011001101010;
      patterns[4409] = 50'b01_0011101101011101_1100101100001101_0111000001010000;
      patterns[4410] = 50'b10_0011101101011101_1100101100001101_0000101100001101;
      patterns[4411] = 50'b11_0011101101011101_1100101100001101_1111101101011101;
      patterns[4412] = 50'b00_0110100010111100_1111101011001011_0110001110000111;
      patterns[4413] = 50'b01_0110100010111100_1111101011001011_0110110111110001;
      patterns[4414] = 50'b10_0110100010111100_1111101011001011_0110100010001000;
      patterns[4415] = 50'b11_0110100010111100_1111101011001011_1111101011111111;
      patterns[4416] = 50'b00_1111110011010111_1010011001001011_1010001100100010;
      patterns[4417] = 50'b01_1111110011010111_1010011001001011_0101011010001100;
      patterns[4418] = 50'b10_1111110011010111_1010011001001011_1010010001000011;
      patterns[4419] = 50'b11_1111110011010111_1010011001001011_1111111011011111;
      patterns[4420] = 50'b00_1010100010000010_0110001110011100_0000110000011110;
      patterns[4421] = 50'b01_1010100010000010_0110001110011100_0100010011100110;
      patterns[4422] = 50'b10_1010100010000010_0110001110011100_0010000010000000;
      patterns[4423] = 50'b11_1010100010000010_0110001110011100_1110101110011110;
      patterns[4424] = 50'b00_1011010000101110_0011110111000011_1111000111110001;
      patterns[4425] = 50'b01_1011010000101110_0011110111000011_0111011001101011;
      patterns[4426] = 50'b10_1011010000101110_0011110111000011_0011010000000010;
      patterns[4427] = 50'b11_1011010000101110_0011110111000011_1011110111101111;
      patterns[4428] = 50'b00_1110001000000110_0011000101110000_0001001101110110;
      patterns[4429] = 50'b01_1110001000000110_0011000101110000_1011000010010110;
      patterns[4430] = 50'b10_1110001000000110_0011000101110000_0010000000000000;
      patterns[4431] = 50'b11_1110001000000110_0011000101110000_1111001101110110;
      patterns[4432] = 50'b00_1010010001010110_0100111111011001_1111010000101111;
      patterns[4433] = 50'b01_1010010001010110_0100111111011001_0101010001111101;
      patterns[4434] = 50'b10_1010010001010110_0100111111011001_0000010001010000;
      patterns[4435] = 50'b11_1010010001010110_0100111111011001_1110111111011111;
      patterns[4436] = 50'b00_0010011111010110_1111111111100011_0010011110111001;
      patterns[4437] = 50'b01_0010011111010110_1111111111100011_0010011111110011;
      patterns[4438] = 50'b10_0010011111010110_1111111111100011_0010011111000010;
      patterns[4439] = 50'b11_0010011111010110_1111111111100011_1111111111110111;
      patterns[4440] = 50'b00_1100000101011001_1111010110111011_1011011100010100;
      patterns[4441] = 50'b01_1100000101011001_1111010110111011_1100101110011110;
      patterns[4442] = 50'b10_1100000101011001_1111010110111011_1100000100011001;
      patterns[4443] = 50'b11_1100000101011001_1111010110111011_1111010111111011;
      patterns[4444] = 50'b00_0110000001110001_0011101101010111_1001101111001000;
      patterns[4445] = 50'b01_0110000001110001_0011101101010111_0010010100011010;
      patterns[4446] = 50'b10_0110000001110001_0011101101010111_0010000001010001;
      patterns[4447] = 50'b11_0110000001110001_0011101101010111_0111101101110111;
      patterns[4448] = 50'b00_0100100111111000_0111100000011010_1100001000010010;
      patterns[4449] = 50'b01_0100100111111000_0111100000011010_1101000111011110;
      patterns[4450] = 50'b10_0100100111111000_0111100000011010_0100100000011000;
      patterns[4451] = 50'b11_0100100111111000_0111100000011010_0111100111111010;
      patterns[4452] = 50'b00_1010111101001110_1010111001000001_0101110110001111;
      patterns[4453] = 50'b01_1010111101001110_1010111001000001_0000000100001101;
      patterns[4454] = 50'b10_1010111101001110_1010111001000001_1010111001000000;
      patterns[4455] = 50'b11_1010111101001110_1010111001000001_1010111101001111;
      patterns[4456] = 50'b00_1010111100000110_1111100100100111_1010100000101101;
      patterns[4457] = 50'b01_1010111100000110_1111100100100111_1011010111011111;
      patterns[4458] = 50'b10_1010111100000110_1111100100100111_1010100100000110;
      patterns[4459] = 50'b11_1010111100000110_1111100100100111_1111111100100111;
      patterns[4460] = 50'b00_1111001001100001_1100001100011000_1011010101111001;
      patterns[4461] = 50'b01_1111001001100001_1100001100011000_0010111101001001;
      patterns[4462] = 50'b10_1111001001100001_1100001100011000_1100001000000000;
      patterns[4463] = 50'b11_1111001001100001_1100001100011000_1111001101111001;
      patterns[4464] = 50'b00_1100111001100011_0010101101011100_1111100110111111;
      patterns[4465] = 50'b01_1100111001100011_0010101101011100_1010001100000111;
      patterns[4466] = 50'b10_1100111001100011_0010101101011100_0000101001000000;
      patterns[4467] = 50'b11_1100111001100011_0010101101011100_1110111101111111;
      patterns[4468] = 50'b00_0111111111000110_0110000100001011_1110000011010001;
      patterns[4469] = 50'b01_0111111111000110_0110000100001011_0001111010111011;
      patterns[4470] = 50'b10_0111111111000110_0110000100001011_0110000100000010;
      patterns[4471] = 50'b11_0111111111000110_0110000100001011_0111111111001111;
      patterns[4472] = 50'b00_1000110011101011_1111001111011000_1000000011000011;
      patterns[4473] = 50'b01_1000110011101011_1111001111011000_1001100100010011;
      patterns[4474] = 50'b10_1000110011101011_1111001111011000_1000000011001000;
      patterns[4475] = 50'b11_1000110011101011_1111001111011000_1111111111111011;
      patterns[4476] = 50'b00_0110100001100100_0010010011101011_1000110101001111;
      patterns[4477] = 50'b01_0110100001100100_0010010011101011_0100001101111001;
      patterns[4478] = 50'b10_0110100001100100_0010010011101011_0010000001100000;
      patterns[4479] = 50'b11_0110100001100100_0010010011101011_0110110011101111;
      patterns[4480] = 50'b00_0100011110111001_0010011001100011_0110111000011100;
      patterns[4481] = 50'b01_0100011110111001_0010011001100011_0010000101010110;
      patterns[4482] = 50'b10_0100011110111001_0010011001100011_0000011000100001;
      patterns[4483] = 50'b11_0100011110111001_0010011001100011_0110011111111011;
      patterns[4484] = 50'b00_1000010110101100_1011101011110011_0100000010011111;
      patterns[4485] = 50'b01_1000010110101100_1011101011110011_1100101010111001;
      patterns[4486] = 50'b10_1000010110101100_1011101011110011_1000000010100000;
      patterns[4487] = 50'b11_1000010110101100_1011101011110011_1011111111111111;
      patterns[4488] = 50'b00_0110101010001101_1000000001010111_1110101011100100;
      patterns[4489] = 50'b01_0110101010001101_1000000001010111_1110101000110110;
      patterns[4490] = 50'b10_0110101010001101_1000000001010111_0000000000000101;
      patterns[4491] = 50'b11_0110101010001101_1000000001010111_1110101011011111;
      patterns[4492] = 50'b00_1000000110111110_0100100101011001_1100101100010111;
      patterns[4493] = 50'b01_1000000110111110_0100100101011001_0011100001100101;
      patterns[4494] = 50'b10_1000000110111110_0100100101011001_0000000100011000;
      patterns[4495] = 50'b11_1000000110111110_0100100101011001_1100100111111111;
      patterns[4496] = 50'b00_1011011001000001_1010011100000000_0101110101000001;
      patterns[4497] = 50'b01_1011011001000001_1010011100000000_0000111101000001;
      patterns[4498] = 50'b10_1011011001000001_1010011100000000_1010011000000000;
      patterns[4499] = 50'b11_1011011001000001_1010011100000000_1011011101000001;
      patterns[4500] = 50'b00_1101101010011110_0010111011001110_0000100101101100;
      patterns[4501] = 50'b01_1101101010011110_0010111011001110_1010101111010000;
      patterns[4502] = 50'b10_1101101010011110_0010111011001110_0000101010001110;
      patterns[4503] = 50'b11_1101101010011110_0010111011001110_1111111011011110;
      patterns[4504] = 50'b00_0110011110010010_0011010100111100_1001110011001110;
      patterns[4505] = 50'b01_0110011110010010_0011010100111100_0011001001010110;
      patterns[4506] = 50'b10_0110011110010010_0011010100111100_0010010100010000;
      patterns[4507] = 50'b11_0110011110010010_0011010100111100_0111011110111110;
      patterns[4508] = 50'b00_1001101001001101_1101001101100000_0110110110101101;
      patterns[4509] = 50'b01_1001101001001101_1101001101100000_1100011011101101;
      patterns[4510] = 50'b10_1001101001001101_1101001101100000_1001001001000000;
      patterns[4511] = 50'b11_1001101001001101_1101001101100000_1101101101101101;
      patterns[4512] = 50'b00_0111101110101001_1101001101100000_0100111100001001;
      patterns[4513] = 50'b01_0111101110101001_1101001101100000_1010100001001001;
      patterns[4514] = 50'b10_0111101110101001_1101001101100000_0101001100100000;
      patterns[4515] = 50'b11_0111101110101001_1101001101100000_1111101111101001;
      patterns[4516] = 50'b00_0001111011010111_1110110101011000_0000110000101111;
      patterns[4517] = 50'b01_0001111011010111_1110110101011000_0011000101111111;
      patterns[4518] = 50'b10_0001111011010111_1110110101011000_0000110001010000;
      patterns[4519] = 50'b11_0001111011010111_1110110101011000_1111111111011111;
      patterns[4520] = 50'b00_1100010100110000_1110101110110011_1011000011100011;
      patterns[4521] = 50'b01_1100010100110000_1110101110110011_1101100101111101;
      patterns[4522] = 50'b10_1100010100110000_1110101110110011_1100000100110000;
      patterns[4523] = 50'b11_1100010100110000_1110101110110011_1110111110110011;
      patterns[4524] = 50'b00_1101011011000011_0110011100010011_0011110111010110;
      patterns[4525] = 50'b01_1101011011000011_0110011100010011_0110111110110000;
      patterns[4526] = 50'b10_1101011011000011_0110011100010011_0100011000000011;
      patterns[4527] = 50'b11_1101011011000011_0110011100010011_1111011111010011;
      patterns[4528] = 50'b00_0110000111011001_1100110100000111_0010111011100000;
      patterns[4529] = 50'b01_0110000111011001_1100110100000111_1001010011010010;
      patterns[4530] = 50'b10_0110000111011001_1100110100000111_0100000100000001;
      patterns[4531] = 50'b11_0110000111011001_1100110100000111_1110110111011111;
      patterns[4532] = 50'b00_0100011101101100_0000010111101011_0100110101010111;
      patterns[4533] = 50'b01_0100011101101100_0000010111101011_0100000110000001;
      patterns[4534] = 50'b10_0100011101101100_0000010111101011_0000010101101000;
      patterns[4535] = 50'b11_0100011101101100_0000010111101011_0100011111101111;
      patterns[4536] = 50'b00_0110010110100110_1111010000110100_0101100111011010;
      patterns[4537] = 50'b01_0110010110100110_1111010000110100_0111000101110010;
      patterns[4538] = 50'b10_0110010110100110_1111010000110100_0110010000100100;
      patterns[4539] = 50'b11_0110010110100110_1111010000110100_1111010110110110;
      patterns[4540] = 50'b00_0000110000101011_0000110110101001_0001100111010100;
      patterns[4541] = 50'b01_0000110000101011_0000110110101001_1111111010000010;
      patterns[4542] = 50'b10_0000110000101011_0000110110101001_0000110000101001;
      patterns[4543] = 50'b11_0000110000101011_0000110110101001_0000110110101011;
      patterns[4544] = 50'b00_0011111001011001_1100010010001001_0000001011100010;
      patterns[4545] = 50'b01_0011111001011001_1100010010001001_0111100111010000;
      patterns[4546] = 50'b10_0011111001011001_1100010010001001_0000010000001001;
      patterns[4547] = 50'b11_0011111001011001_1100010010001001_1111111011011001;
      patterns[4548] = 50'b00_1011111001100011_0101111100100100_0001110110000111;
      patterns[4549] = 50'b01_1011111001100011_0101111100100100_0101111100111111;
      patterns[4550] = 50'b10_1011111001100011_0101111100100100_0001111000100000;
      patterns[4551] = 50'b11_1011111001100011_0101111100100100_1111111101100111;
      patterns[4552] = 50'b00_0110011011010011_0010111001110100_1001010101000111;
      patterns[4553] = 50'b01_0110011011010011_0010111001110100_0011100001011111;
      patterns[4554] = 50'b10_0110011011010011_0010111001110100_0010011001010000;
      patterns[4555] = 50'b11_0110011011010011_0010111001110100_0110111011110111;
      patterns[4556] = 50'b00_1101111111001100_1111101111111011_1101101111000111;
      patterns[4557] = 50'b01_1101111111001100_1111101111111011_1110001111010001;
      patterns[4558] = 50'b10_1101111111001100_1111101111111011_1101101111001000;
      patterns[4559] = 50'b11_1101111111001100_1111101111111011_1111111111111111;
      patterns[4560] = 50'b00_0111111101010010_1010001011110001_0010001001000011;
      patterns[4561] = 50'b01_0111111101010010_1010001011110001_1101110001100001;
      patterns[4562] = 50'b10_0111111101010010_1010001011110001_0010001001010000;
      patterns[4563] = 50'b11_0111111101010010_1010001011110001_1111111111110011;
      patterns[4564] = 50'b00_1111000110011100_0110110010000110_0101111000100010;
      patterns[4565] = 50'b01_1111000110011100_0110110010000110_1000010100010110;
      patterns[4566] = 50'b10_1111000110011100_0110110010000110_0110000010000100;
      patterns[4567] = 50'b11_1111000110011100_0110110010000110_1111110110011110;
      patterns[4568] = 50'b00_1100010011010111_0011100110000110_1111111001011101;
      patterns[4569] = 50'b01_1100010011010111_0011100110000110_1000101101010001;
      patterns[4570] = 50'b10_1100010011010111_0011100110000110_0000000010000110;
      patterns[4571] = 50'b11_1100010011010111_0011100110000110_1111110111010111;
      patterns[4572] = 50'b00_1101110001011010_0100000010000010_0001110011011100;
      patterns[4573] = 50'b01_1101110001011010_0100000010000010_1001101111011000;
      patterns[4574] = 50'b10_1101110001011010_0100000010000010_0100000000000010;
      patterns[4575] = 50'b11_1101110001011010_0100000010000010_1101110011011010;
      patterns[4576] = 50'b00_0010111100010111_0001110111011100_0100110011110011;
      patterns[4577] = 50'b01_0010111100010111_0001110111011100_0001000100111011;
      patterns[4578] = 50'b10_0010111100010111_0001110111011100_0000110100010100;
      patterns[4579] = 50'b11_0010111100010111_0001110111011100_0011111111011111;
      patterns[4580] = 50'b00_1010110110001101_1100011000000110_0111001110010011;
      patterns[4581] = 50'b01_1010110110001101_1100011000000110_1110011110000111;
      patterns[4582] = 50'b10_1010110110001101_1100011000000110_1000010000000100;
      patterns[4583] = 50'b11_1010110110001101_1100011000000110_1110111110001111;
      patterns[4584] = 50'b00_0011000111001110_0011000100110011_0110001100000001;
      patterns[4585] = 50'b01_0011000111001110_0011000100110011_0000000010011011;
      patterns[4586] = 50'b10_0011000111001110_0011000100110011_0011000100000010;
      patterns[4587] = 50'b11_0011000111001110_0011000100110011_0011000111111111;
      patterns[4588] = 50'b00_0111100101111111_0001110110111111_1001011100111110;
      patterns[4589] = 50'b01_0111100101111111_0001110110111111_0101101111000000;
      patterns[4590] = 50'b10_0111100101111111_0001110110111111_0001100100111111;
      patterns[4591] = 50'b11_0111100101111111_0001110110111111_0111110111111111;
      patterns[4592] = 50'b00_0011101101001111_0100101101001011_1000011010011010;
      patterns[4593] = 50'b01_0011101101001111_0100101101001011_1111000000000100;
      patterns[4594] = 50'b10_0011101101001111_0100101101001011_0000101101001011;
      patterns[4595] = 50'b11_0011101101001111_0100101101001011_0111101101001111;
      patterns[4596] = 50'b00_1110000011010100_0000011010010011_1110011101100111;
      patterns[4597] = 50'b01_1110000011010100_0000011010010011_1101101001000001;
      patterns[4598] = 50'b10_1110000011010100_0000011010010011_0000000010010000;
      patterns[4599] = 50'b11_1110000011010100_0000011010010011_1110011011010111;
      patterns[4600] = 50'b00_1000111110100010_1010110110000000_0011110100100010;
      patterns[4601] = 50'b01_1000111110100010_1010110110000000_1110001000100010;
      patterns[4602] = 50'b10_1000111110100010_1010110110000000_1000110110000000;
      patterns[4603] = 50'b11_1000111110100010_1010110110000000_1010111110100010;
      patterns[4604] = 50'b00_0101001010110001_0001011000011010_0110100011001011;
      patterns[4605] = 50'b01_0101001010110001_0001011000011010_0011110010010111;
      patterns[4606] = 50'b10_0101001010110001_0001011000011010_0001001000010000;
      patterns[4607] = 50'b11_0101001010110001_0001011000011010_0101011010111011;
      patterns[4608] = 50'b00_0000110010100111_0000101000100110_0001011011001101;
      patterns[4609] = 50'b01_0000110010100111_0000101000100110_0000001010000001;
      patterns[4610] = 50'b10_0000110010100111_0000101000100110_0000100000100110;
      patterns[4611] = 50'b11_0000110010100111_0000101000100110_0000111010100111;
      patterns[4612] = 50'b00_1010010110011100_1001011010001111_0011110000101011;
      patterns[4613] = 50'b01_1010010110011100_1001011010001111_0000111100001101;
      patterns[4614] = 50'b10_1010010110011100_1001011010001111_1000010010001100;
      patterns[4615] = 50'b11_1010010110011100_1001011010001111_1011011110011111;
      patterns[4616] = 50'b00_1011100011100111_1111100101110010_1011001001011001;
      patterns[4617] = 50'b01_1011100011100111_1111100101110010_1011111101110101;
      patterns[4618] = 50'b10_1011100011100111_1111100101110010_1011100001100010;
      patterns[4619] = 50'b11_1011100011100111_1111100101110010_1111100111110111;
      patterns[4620] = 50'b00_0000101001101000_1110111000110101_1111100010011101;
      patterns[4621] = 50'b01_0000101001101000_1110111000110101_0001110000110011;
      patterns[4622] = 50'b10_0000101001101000_1110111000110101_0000101000100000;
      patterns[4623] = 50'b11_0000101001101000_1110111000110101_1110111001111101;
      patterns[4624] = 50'b00_1011110000100011_1101010001110110_1001000010011001;
      patterns[4625] = 50'b01_1011110000100011_1101010001110110_1110011110101101;
      patterns[4626] = 50'b10_1011110000100011_1101010001110110_1001010000100010;
      patterns[4627] = 50'b11_1011110000100011_1101010001110110_1111110001110111;
      patterns[4628] = 50'b00_1010110111010010_0100011100111101_1111010100001111;
      patterns[4629] = 50'b01_1010110111010010_0100011100111101_0110011010010101;
      patterns[4630] = 50'b10_1010110111010010_0100011100111101_0000010100010000;
      patterns[4631] = 50'b11_1010110111010010_0100011100111101_1110111111111111;
      patterns[4632] = 50'b00_1000010111010010_1011010111111100_0011101111001110;
      patterns[4633] = 50'b01_1000010111010010_1011010111111100_1100111111010110;
      patterns[4634] = 50'b10_1000010111010010_1011010111111100_1000010111010000;
      patterns[4635] = 50'b11_1000010111010010_1011010111111100_1011010111111110;
      patterns[4636] = 50'b00_1001011010011001_0010101010110111_1100000101010000;
      patterns[4637] = 50'b01_1001011010011001_0010101010110111_0110101111100010;
      patterns[4638] = 50'b10_1001011010011001_0010101010110111_0000001010010001;
      patterns[4639] = 50'b11_1001011010011001_0010101010110111_1011111010111111;
      patterns[4640] = 50'b00_0111001011111100_1101000001001111_0100001101001011;
      patterns[4641] = 50'b01_0111001011111100_1101000001001111_1010001010101101;
      patterns[4642] = 50'b10_0111001011111100_1101000001001111_0101000001001100;
      patterns[4643] = 50'b11_0111001011111100_1101000001001111_1111001011111111;
      patterns[4644] = 50'b00_0110111100111000_1110010000100000_0101001101011000;
      patterns[4645] = 50'b01_0110111100111000_1110010000100000_1000101100011000;
      patterns[4646] = 50'b10_0110111100111000_1110010000100000_0110010000100000;
      patterns[4647] = 50'b11_0110111100111000_1110010000100000_1110111100111000;
      patterns[4648] = 50'b00_0011101001000110_0101111000101010_1001100001110000;
      patterns[4649] = 50'b01_0011101001000110_0101111000101010_1101110000011100;
      patterns[4650] = 50'b10_0011101001000110_0101111000101010_0001101000000010;
      patterns[4651] = 50'b11_0011101001000110_0101111000101010_0111111001101110;
      patterns[4652] = 50'b00_1111001110010011_1100111010000010_1100001000010101;
      patterns[4653] = 50'b01_1111001110010011_1100111010000010_0010010100010001;
      patterns[4654] = 50'b10_1111001110010011_1100111010000010_1100001010000010;
      patterns[4655] = 50'b11_1111001110010011_1100111010000010_1111111110010011;
      patterns[4656] = 50'b00_1100001000010001_0011010001110011_1111011010000100;
      patterns[4657] = 50'b01_1100001000010001_0011010001110011_1000110110011110;
      patterns[4658] = 50'b10_1100001000010001_0011010001110011_0000000000010001;
      patterns[4659] = 50'b11_1100001000010001_0011010001110011_1111011001110011;
      patterns[4660] = 50'b00_1010110000111111_0001111101010010_1100101110010001;
      patterns[4661] = 50'b01_1010110000111111_0001111101010010_1000110011101101;
      patterns[4662] = 50'b10_1010110000111111_0001111101010010_0000110000010010;
      patterns[4663] = 50'b11_1010110000111111_0001111101010010_1011111101111111;
      patterns[4664] = 50'b00_1100100111110001_0110000101110100_0010101101100101;
      patterns[4665] = 50'b01_1100100111110001_0110000101110100_0110100001111101;
      patterns[4666] = 50'b10_1100100111110001_0110000101110100_0100000101110000;
      patterns[4667] = 50'b11_1100100111110001_0110000101110100_1110100111110101;
      patterns[4668] = 50'b00_0111101000101000_0101111001101000_1101100010010000;
      patterns[4669] = 50'b01_0111101000101000_0101111001101000_0001101111000000;
      patterns[4670] = 50'b10_0111101000101000_0101111001101000_0101101000101000;
      patterns[4671] = 50'b11_0111101000101000_0101111001101000_0111111001101000;
      patterns[4672] = 50'b00_1111110111110101_0101010110100101_0101001110011010;
      patterns[4673] = 50'b01_1111110111110101_0101010110100101_1010100001010000;
      patterns[4674] = 50'b10_1111110111110101_0101010110100101_0101010110100101;
      patterns[4675] = 50'b11_1111110111110101_0101010110100101_1111110111110101;
      patterns[4676] = 50'b00_0011011011000100_0111110111001111_1011010010010011;
      patterns[4677] = 50'b01_0011011011000100_0111110111001111_1011100011110101;
      patterns[4678] = 50'b10_0011011011000100_0111110111001111_0011010011000100;
      patterns[4679] = 50'b11_0011011011000100_0111110111001111_0111111111001111;
      patterns[4680] = 50'b00_1001111101111010_1100100101010100_0110100011001110;
      patterns[4681] = 50'b01_1001111101111010_1100100101010100_1101011000100110;
      patterns[4682] = 50'b10_1001111101111010_1100100101010100_1000100101010000;
      patterns[4683] = 50'b11_1001111101111010_1100100101010100_1101111101111110;
      patterns[4684] = 50'b00_0101011000101000_0110111101000111_1100010101101111;
      patterns[4685] = 50'b01_0101011000101000_0110111101000111_1110011011100001;
      patterns[4686] = 50'b10_0101011000101000_0110111101000111_0100011000000000;
      patterns[4687] = 50'b11_0101011000101000_0110111101000111_0111111101101111;
      patterns[4688] = 50'b00_1110110010000011_1111000110101111_1101111000110010;
      patterns[4689] = 50'b01_1110110010000011_1111000110101111_1111101011010100;
      patterns[4690] = 50'b10_1110110010000011_1111000110101111_1110000010000011;
      patterns[4691] = 50'b11_1110110010000011_1111000110101111_1111110110101111;
      patterns[4692] = 50'b00_0000100110001111_0010100010101101_0011001000111100;
      patterns[4693] = 50'b01_0000100110001111_0010100010101101_1110000011100010;
      patterns[4694] = 50'b10_0000100110001111_0010100010101101_0000100010001101;
      patterns[4695] = 50'b11_0000100110001111_0010100010101101_0010100110101111;
      patterns[4696] = 50'b00_1101001111001011_1001111100000010_0111001011001101;
      patterns[4697] = 50'b01_1101001111001011_1001111100000010_0011010011001001;
      patterns[4698] = 50'b10_1101001111001011_1001111100000010_1001001100000010;
      patterns[4699] = 50'b11_1101001111001011_1001111100000010_1101111111001011;
      patterns[4700] = 50'b00_1101101000111010_0100001110101001_0001110111100011;
      patterns[4701] = 50'b01_1101101000111010_0100001110101001_1001011010010001;
      patterns[4702] = 50'b10_1101101000111010_0100001110101001_0100001000101000;
      patterns[4703] = 50'b11_1101101000111010_0100001110101001_1101101110111011;
      patterns[4704] = 50'b00_0101000100010100_1000110100100011_1101111000110111;
      patterns[4705] = 50'b01_0101000100010100_1000110100100011_1100001111110001;
      patterns[4706] = 50'b10_0101000100010100_1000110100100011_0000000100000000;
      patterns[4707] = 50'b11_0101000100010100_1000110100100011_1101110100110111;
      patterns[4708] = 50'b00_0001010110111001_1100100001010101_1101111000001110;
      patterns[4709] = 50'b01_0001010110111001_1100100001010101_0100110101100100;
      patterns[4710] = 50'b10_0001010110111001_1100100001010101_0000000000010001;
      patterns[4711] = 50'b11_0001010110111001_1100100001010101_1101110111111101;
      patterns[4712] = 50'b00_0000001001101000_1000011001101111_1000100011010111;
      patterns[4713] = 50'b01_0000001001101000_1000011001101111_0111101111111001;
      patterns[4714] = 50'b10_0000001001101000_1000011001101111_0000001001101000;
      patterns[4715] = 50'b11_0000001001101000_1000011001101111_1000011001101111;
      patterns[4716] = 50'b00_1010111000000000_0011110111000111_1110101111000111;
      patterns[4717] = 50'b01_1010111000000000_0011110111000111_0111000000111001;
      patterns[4718] = 50'b10_1010111000000000_0011110111000111_0010110000000000;
      patterns[4719] = 50'b11_1010111000000000_0011110111000111_1011111111000111;
      patterns[4720] = 50'b00_0010010001000010_1111100011000111_0001110100001001;
      patterns[4721] = 50'b01_0010010001000010_1111100011000111_0010101101111011;
      patterns[4722] = 50'b10_0010010001000010_1111100011000111_0010000001000010;
      patterns[4723] = 50'b11_0010010001000010_1111100011000111_1111110011000111;
      patterns[4724] = 50'b00_0110000011010111_1100111010100001_0010111101111000;
      patterns[4725] = 50'b01_0110000011010111_1100111010100001_1001001000110110;
      patterns[4726] = 50'b10_0110000011010111_1100111010100001_0100000010000001;
      patterns[4727] = 50'b11_0110000011010111_1100111010100001_1110111011110111;
      patterns[4728] = 50'b00_0010011111100001_0100001101101101_0110101101001110;
      patterns[4729] = 50'b01_0010011111100001_0100001101101101_1110010001110100;
      patterns[4730] = 50'b10_0010011111100001_0100001101101101_0000001101100001;
      patterns[4731] = 50'b11_0010011111100001_0100001101101101_0110011111101101;
      patterns[4732] = 50'b00_0001001110001111_0010101100010000_0011111010011111;
      patterns[4733] = 50'b01_0001001110001111_0010101100010000_1110100001111111;
      patterns[4734] = 50'b10_0001001110001111_0010101100010000_0000001100000000;
      patterns[4735] = 50'b11_0001001110001111_0010101100010000_0011101110011111;
      patterns[4736] = 50'b00_1000010000111011_0101001110111100_1101011111110111;
      patterns[4737] = 50'b01_1000010000111011_0101001110111100_0011000001111111;
      patterns[4738] = 50'b10_1000010000111011_0101001110111100_0000000000111000;
      patterns[4739] = 50'b11_1000010000111011_0101001110111100_1101011110111111;
      patterns[4740] = 50'b00_0101000100000001_1101010011111000_0010010111111001;
      patterns[4741] = 50'b01_0101000100000001_1101010011111000_0111110000001001;
      patterns[4742] = 50'b10_0101000100000001_1101010011111000_0101000000000000;
      patterns[4743] = 50'b11_0101000100000001_1101010011111000_1101010111111001;
      patterns[4744] = 50'b00_0011011101001101_0001111000001111_0101010101011100;
      patterns[4745] = 50'b01_0011011101001101_0001111000001111_0001100100111110;
      patterns[4746] = 50'b10_0011011101001101_0001111000001111_0001011000001101;
      patterns[4747] = 50'b11_0011011101001101_0001111000001111_0011111101001111;
      patterns[4748] = 50'b00_1100000101000100_1010111000010101_0110111101011001;
      patterns[4749] = 50'b01_1100000101000100_1010111000010101_0001001100101111;
      patterns[4750] = 50'b10_1100000101000100_1010111000010101_1000000000000100;
      patterns[4751] = 50'b11_1100000101000100_1010111000010101_1110111101010101;
      patterns[4752] = 50'b00_1010101010110101_0001111101010111_1100101000001100;
      patterns[4753] = 50'b01_1010101010110101_0001111101010111_1000101101011110;
      patterns[4754] = 50'b10_1010101010110101_0001111101010111_0000101000010101;
      patterns[4755] = 50'b11_1010101010110101_0001111101010111_1011111111110111;
      patterns[4756] = 50'b00_0100001110101010_1111001101011110_0011011100001000;
      patterns[4757] = 50'b01_0100001110101010_1111001101011110_0101000001001100;
      patterns[4758] = 50'b10_0100001110101010_1111001101011110_0100001100001010;
      patterns[4759] = 50'b11_0100001110101010_1111001101011110_1111001111111110;
      patterns[4760] = 50'b00_0101001111100111_0101101100111000_1010111100011111;
      patterns[4761] = 50'b01_0101001111100111_0101101100111000_1111100010101111;
      patterns[4762] = 50'b10_0101001111100111_0101101100111000_0101001100100000;
      patterns[4763] = 50'b11_0101001111100111_0101101100111000_0101101111111111;
      patterns[4764] = 50'b00_0000110011100000_0100101111110111_0101100011010111;
      patterns[4765] = 50'b01_0000110011100000_0100101111110111_1100000011101001;
      patterns[4766] = 50'b10_0000110011100000_0100101111110111_0000100011100000;
      patterns[4767] = 50'b11_0000110011100000_0100101111110111_0100111111110111;
      patterns[4768] = 50'b00_0111010101100100_0011100110101000_1010111100001100;
      patterns[4769] = 50'b01_0111010101100100_0011100110101000_0011101110111100;
      patterns[4770] = 50'b10_0111010101100100_0011100110101000_0011000100100000;
      patterns[4771] = 50'b11_0111010101100100_0011100110101000_0111110111101100;
      patterns[4772] = 50'b00_1100110001001101_0011010101110010_0000000110111111;
      patterns[4773] = 50'b01_1100110001001101_0011010101110010_1001011011011011;
      patterns[4774] = 50'b10_1100110001001101_0011010101110010_0000010001000000;
      patterns[4775] = 50'b11_1100110001001101_0011010101110010_1111110101111111;
      patterns[4776] = 50'b00_1101101110110011_0011111001100100_0001101000010111;
      patterns[4777] = 50'b01_1101101110110011_0011111001100100_1001110101001111;
      patterns[4778] = 50'b10_1101101110110011_0011111001100100_0001101000100000;
      patterns[4779] = 50'b11_1101101110110011_0011111001100100_1111111111110111;
      patterns[4780] = 50'b00_0110010100000101_1110001000111100_0100011101000001;
      patterns[4781] = 50'b01_0110010100000101_1110001000111100_1000001011001001;
      patterns[4782] = 50'b10_0110010100000101_1110001000111100_0110000000000100;
      patterns[4783] = 50'b11_0110010100000101_1110001000111100_1110011100111101;
      patterns[4784] = 50'b00_0100111000010110_1101001111000001_0010000111010111;
      patterns[4785] = 50'b01_0100111000010110_1101001111000001_0111101001010101;
      patterns[4786] = 50'b10_0100111000010110_1101001111000001_0100001000000000;
      patterns[4787] = 50'b11_0100111000010110_1101001111000001_1101111111010111;
      patterns[4788] = 50'b00_0011011111110000_1001001001100011_1100101001010011;
      patterns[4789] = 50'b01_0011011111110000_1001001001100011_1010010110001101;
      patterns[4790] = 50'b10_0011011111110000_1001001001100011_0001001001100000;
      patterns[4791] = 50'b11_0011011111110000_1001001001100011_1011011111110011;
      patterns[4792] = 50'b00_1011000000111101_0100100110100100_1111100111100001;
      patterns[4793] = 50'b01_1011000000111101_0100100110100100_0110011010011001;
      patterns[4794] = 50'b10_1011000000111101_0100100110100100_0000000000100100;
      patterns[4795] = 50'b11_1011000000111101_0100100110100100_1111100110111101;
      patterns[4796] = 50'b00_0101010111111100_1000101000100011_1110000000011111;
      patterns[4797] = 50'b01_0101010111111100_1000101000100011_1100101111011001;
      patterns[4798] = 50'b10_0101010111111100_1000101000100011_0000000000100000;
      patterns[4799] = 50'b11_0101010111111100_1000101000100011_1101111111111111;
      patterns[4800] = 50'b00_0111111101011001_1011100010101000_0011100000000001;
      patterns[4801] = 50'b01_0111111101011001_1011100010101000_1100011010110001;
      patterns[4802] = 50'b10_0111111101011001_1011100010101000_0011100000001000;
      patterns[4803] = 50'b11_0111111101011001_1011100010101000_1111111111111001;
      patterns[4804] = 50'b00_0011001001110100_0000110011011101_0011111101010001;
      patterns[4805] = 50'b01_0011001001110100_0000110011011101_0010010110010111;
      patterns[4806] = 50'b10_0011001001110100_0000110011011101_0000000001010100;
      patterns[4807] = 50'b11_0011001001110100_0000110011011101_0011111011111101;
      patterns[4808] = 50'b00_0110101001101100_1011000011000110_0001101100110010;
      patterns[4809] = 50'b01_0110101001101100_1011000011000110_1011100110100110;
      patterns[4810] = 50'b10_0110101001101100_1011000011000110_0010000001000100;
      patterns[4811] = 50'b11_0110101001101100_1011000011000110_1111101011101110;
      patterns[4812] = 50'b00_1001011011010110_0010111001100111_1100010100111101;
      patterns[4813] = 50'b01_1001011011010110_0010111001100111_0110100001101111;
      patterns[4814] = 50'b10_1001011011010110_0010111001100111_0000011001000110;
      patterns[4815] = 50'b11_1001011011010110_0010111001100111_1011111011110111;
      patterns[4816] = 50'b00_0100001010110010_0111100111111100_1011110010101110;
      patterns[4817] = 50'b01_0100001010110010_0111100111111100_1100100010110110;
      patterns[4818] = 50'b10_0100001010110010_0111100111111100_0100000010110000;
      patterns[4819] = 50'b11_0100001010110010_0111100111111100_0111101111111110;
      patterns[4820] = 50'b00_1010101011000010_1101111111100001_1000101010100011;
      patterns[4821] = 50'b01_1010101011000010_1101111111100001_1100101011100001;
      patterns[4822] = 50'b10_1010101011000010_1101111111100001_1000101011000000;
      patterns[4823] = 50'b11_1010101011000010_1101111111100001_1111111111100011;
      patterns[4824] = 50'b00_0110011001101000_0011010011000000_1001101100101000;
      patterns[4825] = 50'b01_0110011001101000_0011010011000000_0011000110101000;
      patterns[4826] = 50'b10_0110011001101000_0011010011000000_0010010001000000;
      patterns[4827] = 50'b11_0110011001101000_0011010011000000_0111011011101000;
      patterns[4828] = 50'b00_1101101111011111_0101100001110011_0011010001010010;
      patterns[4829] = 50'b01_1101101111011111_0101100001110011_1000001101101100;
      patterns[4830] = 50'b10_1101101111011111_0101100001110011_0101100001010011;
      patterns[4831] = 50'b11_1101101111011111_0101100001110011_1101101111111111;
      patterns[4832] = 50'b00_0001010101110011_0101011101010110_0110110011001001;
      patterns[4833] = 50'b01_0001010101110011_0101011101010110_1011111000011101;
      patterns[4834] = 50'b10_0001010101110011_0101011101010110_0001010101010010;
      patterns[4835] = 50'b11_0001010101110011_0101011101010110_0101011101110111;
      patterns[4836] = 50'b00_0101001011001000_1101110110011101_0011000001100101;
      patterns[4837] = 50'b01_0101001011001000_1101110110011101_0111010100101011;
      patterns[4838] = 50'b10_0101001011001000_1101110110011101_0101000010001000;
      patterns[4839] = 50'b11_0101001011001000_1101110110011101_1101111111011101;
      patterns[4840] = 50'b00_1101010010010001_1101110000111110_1011000011001111;
      patterns[4841] = 50'b01_1101010010010001_1101110000111110_1111100001010011;
      patterns[4842] = 50'b10_1101010010010001_1101110000111110_1101010000010000;
      patterns[4843] = 50'b11_1101010010010001_1101110000111110_1101110010111111;
      patterns[4844] = 50'b00_0110101101100101_1111101000010000_0110010101110101;
      patterns[4845] = 50'b01_0110101101100101_1111101000010000_0111000101010101;
      patterns[4846] = 50'b10_0110101101100101_1111101000010000_0110101000000000;
      patterns[4847] = 50'b11_0110101101100101_1111101000010000_1111101101110101;
      patterns[4848] = 50'b00_0010000100011011_1111010101010110_0001011001110001;
      patterns[4849] = 50'b01_0010000100011011_1111010101010110_0010101111000101;
      patterns[4850] = 50'b10_0010000100011011_1111010101010110_0010000100010010;
      patterns[4851] = 50'b11_0010000100011011_1111010101010110_1111010101011111;
      patterns[4852] = 50'b00_0101100001000101_0110010100101010_1011110101101111;
      patterns[4853] = 50'b01_0101100001000101_0110010100101010_1111001100011011;
      patterns[4854] = 50'b10_0101100001000101_0110010100101010_0100000000000000;
      patterns[4855] = 50'b11_0101100001000101_0110010100101010_0111110101101111;
      patterns[4856] = 50'b00_0011110010001110_0011111001110001_0111101011111111;
      patterns[4857] = 50'b01_0011110010001110_0011111001110001_1111111000011101;
      patterns[4858] = 50'b10_0011110010001110_0011111001110001_0011110000000000;
      patterns[4859] = 50'b11_0011110010001110_0011111001110001_0011111011111111;
      patterns[4860] = 50'b00_1011000111010001_0011100010000101_1110101001010110;
      patterns[4861] = 50'b01_1011000111010001_0011100010000101_0111100101001100;
      patterns[4862] = 50'b10_1011000111010001_0011100010000101_0011000010000001;
      patterns[4863] = 50'b11_1011000111010001_0011100010000101_1011100111010101;
      patterns[4864] = 50'b00_1100010001010000_0011100101101011_1111110110111011;
      patterns[4865] = 50'b01_1100010001010000_0011100101101011_1000101011100101;
      patterns[4866] = 50'b10_1100010001010000_0011100101101011_0000000001000000;
      patterns[4867] = 50'b11_1100010001010000_0011100101101011_1111110101111011;
      patterns[4868] = 50'b00_0011001101110101_1001010001001010_1100011110111111;
      patterns[4869] = 50'b01_0011001101110101_1001010001001010_1001111100101011;
      patterns[4870] = 50'b10_0011001101110101_1001010001001010_0001000001000000;
      patterns[4871] = 50'b11_0011001101110101_1001010001001010_1011011101111111;
      patterns[4872] = 50'b00_0001111101110011_0101010100001110_0111010010000001;
      patterns[4873] = 50'b01_0001111101110011_0101010100001110_1100101001100101;
      patterns[4874] = 50'b10_0001111101110011_0101010100001110_0001010100000010;
      patterns[4875] = 50'b11_0001111101110011_0101010100001110_0101111101111111;
      patterns[4876] = 50'b00_0101001000011000_0111111000100110_1101000000111110;
      patterns[4877] = 50'b01_0101001000011000_0111111000100110_1101001111110010;
      patterns[4878] = 50'b10_0101001000011000_0111111000100110_0101001000000000;
      patterns[4879] = 50'b11_0101001000011000_0111111000100110_0111111000111110;
      patterns[4880] = 50'b00_1000100101101001_1101111101000110_0110100010101111;
      patterns[4881] = 50'b01_1000100101101001_1101111101000110_1010101000100011;
      patterns[4882] = 50'b10_1000100101101001_1101111101000110_1000100101000000;
      patterns[4883] = 50'b11_1000100101101001_1101111101000110_1101111101101111;
      patterns[4884] = 50'b00_1010100010000010_1001101000010101_0100001010010111;
      patterns[4885] = 50'b01_1010100010000010_1001101000010101_0000111001101101;
      patterns[4886] = 50'b10_1010100010000010_1001101000010101_1000100000000000;
      patterns[4887] = 50'b11_1010100010000010_1001101000010101_1011101010010111;
      patterns[4888] = 50'b00_1010010111101110_0000101001111100_1011000001101010;
      patterns[4889] = 50'b01_1010010111101110_0000101001111100_1001101101110010;
      patterns[4890] = 50'b10_1010010111101110_0000101001111100_0000000001101100;
      patterns[4891] = 50'b11_1010010111101110_0000101001111100_1010111111111110;
      patterns[4892] = 50'b00_0110111101111100_0101011101100010_1100011011011110;
      patterns[4893] = 50'b01_0110111101111100_0101011101100010_0001100000011010;
      patterns[4894] = 50'b10_0110111101111100_0101011101100010_0100011101100000;
      patterns[4895] = 50'b11_0110111101111100_0101011101100010_0111111101111110;
      patterns[4896] = 50'b00_0001011110001111_1001110100001100_1011010010011011;
      patterns[4897] = 50'b01_0001011110001111_1001110100001100_0111101010000011;
      patterns[4898] = 50'b10_0001011110001111_1001110100001100_0001010100001100;
      patterns[4899] = 50'b11_0001011110001111_1001110100001100_1001111110001111;
      patterns[4900] = 50'b00_0101100011010111_0100111110011000_1010100001101111;
      patterns[4901] = 50'b01_0101100011010111_0100111110011000_0000100100111111;
      patterns[4902] = 50'b10_0101100011010111_0100111110011000_0100100010010000;
      patterns[4903] = 50'b11_0101100011010111_0100111110011000_0101111111011111;
      patterns[4904] = 50'b00_1000011110011100_1111100100111110_1000000011011010;
      patterns[4905] = 50'b01_1000011110011100_1111100100111110_1000111001011110;
      patterns[4906] = 50'b10_1000011110011100_1111100100111110_1000000100011100;
      patterns[4907] = 50'b11_1000011110011100_1111100100111110_1111111110111110;
      patterns[4908] = 50'b00_0010110110100100_1110000000111000_0000110111011100;
      patterns[4909] = 50'b01_0010110110100100_1110000000111000_0100110101101100;
      patterns[4910] = 50'b10_0010110110100100_1110000000111000_0010000000100000;
      patterns[4911] = 50'b11_0010110110100100_1110000000111000_1110110110111100;
      patterns[4912] = 50'b00_1110101101110001_1110101100110001_1101011010100010;
      patterns[4913] = 50'b01_1110101101110001_1110101100110001_0000000001000000;
      patterns[4914] = 50'b10_1110101101110001_1110101100110001_1110101100110001;
      patterns[4915] = 50'b11_1110101101110001_1110101100110001_1110101101110001;
      patterns[4916] = 50'b00_1000000100111110_0111101101101111_1111110010101101;
      patterns[4917] = 50'b01_1000000100111110_0111101101101111_0000010111001111;
      patterns[4918] = 50'b10_1000000100111110_0111101101101111_0000000100101110;
      patterns[4919] = 50'b11_1000000100111110_0111101101101111_1111101101111111;
      patterns[4920] = 50'b00_1001100001011011_0001000110001110_1010100111101001;
      patterns[4921] = 50'b01_1001100001011011_0001000110001110_1000011011001101;
      patterns[4922] = 50'b10_1001100001011011_0001000110001110_0001000000001010;
      patterns[4923] = 50'b11_1001100001011011_0001000110001110_1001100111011111;
      patterns[4924] = 50'b00_1010010000000110_1100011100101011_0110101100110001;
      patterns[4925] = 50'b01_1010010000000110_1100011100101011_1101110011011011;
      patterns[4926] = 50'b10_1010010000000110_1100011100101011_1000010000000010;
      patterns[4927] = 50'b11_1010010000000110_1100011100101011_1110011100101111;
      patterns[4928] = 50'b00_1110010010001010_1100010100010001_1010100110011011;
      patterns[4929] = 50'b01_1110010010001010_1100010100010001_0001111101111001;
      patterns[4930] = 50'b10_1110010010001010_1100010100010001_1100010000000000;
      patterns[4931] = 50'b11_1110010010001010_1100010100010001_1110010110011011;
      patterns[4932] = 50'b00_1100000111010110_0110010101000110_0010011100011100;
      patterns[4933] = 50'b01_1100000111010110_0110010101000110_0101110010010000;
      patterns[4934] = 50'b10_1100000111010110_0110010101000110_0100000101000110;
      patterns[4935] = 50'b11_1100000111010110_0110010101000110_1110010111010110;
      patterns[4936] = 50'b00_1010100011000111_0001101000100110_1100001011101101;
      patterns[4937] = 50'b01_1010100011000111_0001101000100110_1000111010100001;
      patterns[4938] = 50'b10_1010100011000111_0001101000100110_0000100000000110;
      patterns[4939] = 50'b11_1010100011000111_0001101000100110_1011101011100111;
      patterns[4940] = 50'b00_1100000110100111_0010101010100000_1110110001000111;
      patterns[4941] = 50'b01_1100000110100111_0010101010100000_1001011100000111;
      patterns[4942] = 50'b10_1100000110100111_0010101010100000_0000000010100000;
      patterns[4943] = 50'b11_1100000110100111_0010101010100000_1110101110100111;
      patterns[4944] = 50'b00_1111001111111110_1111011100110100_1110101100110010;
      patterns[4945] = 50'b01_1111001111111110_1111011100110100_1111110011001010;
      patterns[4946] = 50'b10_1111001111111110_1111011100110100_1111001100110100;
      patterns[4947] = 50'b11_1111001111111110_1111011100110100_1111011111111110;
      patterns[4948] = 50'b00_0000110011011011_1001111001100000_1010101100111011;
      patterns[4949] = 50'b01_0000110011011011_1001111001100000_0110111001111011;
      patterns[4950] = 50'b10_0000110011011011_1001111001100000_0000110001000000;
      patterns[4951] = 50'b11_0000110011011011_1001111001100000_1001111011111011;
      patterns[4952] = 50'b00_1010011010110110_0100000101001010_1110100000000000;
      patterns[4953] = 50'b01_1010011010110110_0100000101001010_0110010101101100;
      patterns[4954] = 50'b10_1010011010110110_0100000101001010_0000000000000010;
      patterns[4955] = 50'b11_1010011010110110_0100000101001010_1110011111111110;
      patterns[4956] = 50'b00_1101111000101101_1101010110111101_1011001111101010;
      patterns[4957] = 50'b01_1101111000101101_1101010110111101_0000100001110000;
      patterns[4958] = 50'b10_1101111000101101_1101010110111101_1101010000101101;
      patterns[4959] = 50'b11_1101111000101101_1101010110111101_1101111110111101;
      patterns[4960] = 50'b00_0111101000001100_1101000001010000_0100101001011100;
      patterns[4961] = 50'b01_0111101000001100_1101000001010000_1010100110111100;
      patterns[4962] = 50'b10_0111101000001100_1101000001010000_0101000000000000;
      patterns[4963] = 50'b11_0111101000001100_1101000001010000_1111101001011100;
      patterns[4964] = 50'b00_0001100101000001_0010010000000010_0011110101000011;
      patterns[4965] = 50'b01_0001100101000001_0010010000000010_1111010100111111;
      patterns[4966] = 50'b10_0001100101000001_0010010000000010_0000000000000000;
      patterns[4967] = 50'b11_0001100101000001_0010010000000010_0011110101000011;
      patterns[4968] = 50'b00_0010101011011010_0011001011110111_0101110111010001;
      patterns[4969] = 50'b01_0010101011011010_0011001011110111_1111011111100011;
      patterns[4970] = 50'b10_0010101011011010_0011001011110111_0010001011010010;
      patterns[4971] = 50'b11_0010101011011010_0011001011110111_0011101011111111;
      patterns[4972] = 50'b00_1111010101000101_1010000110101100_1001011011110001;
      patterns[4973] = 50'b01_1111010101000101_1010000110101100_0101001110011001;
      patterns[4974] = 50'b10_1111010101000101_1010000110101100_1010000100000100;
      patterns[4975] = 50'b11_1111010101000101_1010000110101100_1111010111101101;
      patterns[4976] = 50'b00_0001111100001110_0100100111110011_0110100100000001;
      patterns[4977] = 50'b01_0001111100001110_0100100111110011_1101010100011011;
      patterns[4978] = 50'b10_0001111100001110_0100100111110011_0000100100000010;
      patterns[4979] = 50'b11_0001111100001110_0100100111110011_0101111111111111;
      patterns[4980] = 50'b00_1111011000101001_0100000011011001_0011011100000010;
      patterns[4981] = 50'b01_1111011000101001_0100000011011001_1011010101010000;
      patterns[4982] = 50'b10_1111011000101001_0100000011011001_0100000000001001;
      patterns[4983] = 50'b11_1111011000101001_0100000011011001_1111011011111001;
      patterns[4984] = 50'b00_1110000001101000_0110100101010001_0100100110111001;
      patterns[4985] = 50'b01_1110000001101000_0110100101010001_0111011100010111;
      patterns[4986] = 50'b10_1110000001101000_0110100101010001_0110000001000000;
      patterns[4987] = 50'b11_1110000001101000_0110100101010001_1110100101111001;
      patterns[4988] = 50'b00_1100100101100000_0000000001100000_1100100111000000;
      patterns[4989] = 50'b01_1100100101100000_0000000001100000_1100100100000000;
      patterns[4990] = 50'b10_1100100101100000_0000000001100000_0000000001100000;
      patterns[4991] = 50'b11_1100100101100000_0000000001100000_1100100101100000;
      patterns[4992] = 50'b00_0011010100010011_1111110111101010_0011001011111101;
      patterns[4993] = 50'b01_0011010100010011_1111110111101010_0011011100101001;
      patterns[4994] = 50'b10_0011010100010011_1111110111101010_0011010100000010;
      patterns[4995] = 50'b11_0011010100010011_1111110111101010_1111110111111011;
      patterns[4996] = 50'b00_1001110000100100_1101001001010101_0110111001111001;
      patterns[4997] = 50'b01_1001110000100100_1101001001010101_1100100111001111;
      patterns[4998] = 50'b10_1001110000100100_1101001001010101_1001000000000100;
      patterns[4999] = 50'b11_1001110000100100_1101001001010101_1101111001110101;
      patterns[5000] = 50'b00_0111001111011110_1010110001000010_0010000000100000;
      patterns[5001] = 50'b01_0111001111011110_1010110001000010_1100011110011100;
      patterns[5002] = 50'b10_0111001111011110_1010110001000010_0010000001000010;
      patterns[5003] = 50'b11_0111001111011110_1010110001000010_1111111111011110;
      patterns[5004] = 50'b00_0110101010111111_1111010111000111_0110000010000110;
      patterns[5005] = 50'b01_0110101010111111_1111010111000111_0111010011111000;
      patterns[5006] = 50'b10_0110101010111111_1111010111000111_0110000010000111;
      patterns[5007] = 50'b11_0110101010111111_1111010111000111_1111111111111111;
      patterns[5008] = 50'b00_1110111100001001_0111110101011100_0110110001100101;
      patterns[5009] = 50'b01_1110111100001001_0111110101011100_0111000110101101;
      patterns[5010] = 50'b10_1110111100001001_0111110101011100_0110110100001000;
      patterns[5011] = 50'b11_1110111100001001_0111110101011100_1111111101011101;
      patterns[5012] = 50'b00_1001100101001001_1101011011111000_0111000001000001;
      patterns[5013] = 50'b01_1001100101001001_1101011011111000_1100001001010001;
      patterns[5014] = 50'b10_1001100101001001_1101011011111000_1001000001001000;
      patterns[5015] = 50'b11_1001100101001001_1101011011111000_1101111111111001;
      patterns[5016] = 50'b00_1111010111011010_1111010101001011_1110101100100101;
      patterns[5017] = 50'b01_1111010111011010_1111010101001011_0000000010001111;
      patterns[5018] = 50'b10_1111010111011010_1111010101001011_1111010101001010;
      patterns[5019] = 50'b11_1111010111011010_1111010101001011_1111010111011011;
      patterns[5020] = 50'b00_1101111111011001_0000010001101111_1110010001001000;
      patterns[5021] = 50'b01_1101111111011001_0000010001101111_1101101101101010;
      patterns[5022] = 50'b10_1101111111011001_0000010001101111_0000010001001001;
      patterns[5023] = 50'b11_1101111111011001_0000010001101111_1101111111111111;

      for (i = 0; i < 5024; i = i + 1)
      begin
        ALUOP = patterns[i][49:48];
        A = patterns[i][47:32];
        B = patterns[i][31:16];
        #10;
        if (patterns[i][15:0] !== 16'hx)
        begin
          if (RESULT !== patterns[i][15:0])
          begin
            $display("%d:RESULT: (assertion error). Expected %h, found %h", i, patterns[i][15:0], RESULT);
            $finish;
          end
        end
      end

      $display("All tests passed.");
    end
    endmodule
