--  A testbench for alu_RESULT_tb
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

entity alu_RESULT_tb is
end alu_RESULT_tb;

architecture behav of alu_RESULT_tb is
  component main
    port (
      A: in std_logic_vector(15 downto 0); -- First input to ALU
      B: in std_logic_vector(15 downto 0); -- Second input to ALU
      ALUOP: in std_logic_vector(1 downto 0); -- Operation selection input
      RESULT: out std_logic_vector(15 downto 0); -- The result of this ALU operation
      FLAG: out std_logic_vector(3 downto 0) -- The flags associated with the result of this ALU operation
                                             -- 
                                             -- 0. Z (zero)
                                             -- 1. N (negative)
                                             -- 2. C (carry)
                                             -- 3. V (overflow)
      );
  end component;

  signal A : std_logic_vector(15 downto 0);
  signal B : std_logic_vector(15 downto 0);
  signal ALUOP : std_logic_vector(1 downto 0);
  signal RESULT : std_logic_vector(15 downto 0);
  signal FLAG : std_logic_vector(3 downto 0);
  function to_string ( a: std_logic_vector) return string is
      variable b : string (1 to a'length) := (others => NUL);
      variable stri : integer := 1; 
  begin
      for i in a'range loop
          b(stri) := std_logic'image(a((i)))(2);
      stri := stri+1;
      end loop;
      return b;
  end function;
begin
  main_0 : main port map (
    A => A,
    B => B,
    ALUOP => ALUOP,
    RESULT => RESULT,
    FLAG => FLAG );
  process
    type pattern_type is record
      ALUOP : std_logic_vector(1 downto 0);
      A : std_logic_vector(15 downto 0);
      B : std_logic_vector(15 downto 0);
      RESULT : std_logic_vector(15 downto 0);
    end record;
    type pattern_array is array (natural range <>) of pattern_type;
    constant patterns : pattern_array := (
      ("00", "0000000000000000", "0000000000000000", "0000000000000000"), -- i=0
      ("01", "0000000000000000", "0000000000000000", "0000000000000000"), -- i=1
      ("10", "0000000000000000", "0000000000000000", "0000000000000000"), -- i=2
      ("11", "0000000000000000", "0000000000000000", "0000000000000000"), -- i=3
      ("00", "0000000000000000", "0000000000000001", "0000000000000001"), -- i=4
      ("01", "0000000000000000", "0000000000000001", "1111111111111111"), -- i=5
      ("10", "0000000000000000", "0000000000000001", "0000000000000000"), -- i=6
      ("11", "0000000000000000", "0000000000000001", "0000000000000001"), -- i=7
      ("00", "0000000000000000", "0000000000000010", "0000000000000010"), -- i=8
      ("01", "0000000000000000", "0000000000000010", "1111111111111110"), -- i=9
      ("10", "0000000000000000", "0000000000000010", "0000000000000000"), -- i=10
      ("11", "0000000000000000", "0000000000000010", "0000000000000010"), -- i=11
      ("00", "0000000000000000", "0000000000000011", "0000000000000011"), -- i=12
      ("01", "0000000000000000", "0000000000000011", "1111111111111101"), -- i=13
      ("10", "0000000000000000", "0000000000000011", "0000000000000000"), -- i=14
      ("11", "0000000000000000", "0000000000000011", "0000000000000011"), -- i=15
      ("00", "0000000000000000", "0000000000000100", "0000000000000100"), -- i=16
      ("01", "0000000000000000", "0000000000000100", "1111111111111100"), -- i=17
      ("10", "0000000000000000", "0000000000000100", "0000000000000000"), -- i=18
      ("11", "0000000000000000", "0000000000000100", "0000000000000100"), -- i=19
      ("00", "0000000000000000", "0000000000000101", "0000000000000101"), -- i=20
      ("01", "0000000000000000", "0000000000000101", "1111111111111011"), -- i=21
      ("10", "0000000000000000", "0000000000000101", "0000000000000000"), -- i=22
      ("11", "0000000000000000", "0000000000000101", "0000000000000101"), -- i=23
      ("00", "0000000000000000", "0000000000000110", "0000000000000110"), -- i=24
      ("01", "0000000000000000", "0000000000000110", "1111111111111010"), -- i=25
      ("10", "0000000000000000", "0000000000000110", "0000000000000000"), -- i=26
      ("11", "0000000000000000", "0000000000000110", "0000000000000110"), -- i=27
      ("00", "0000000000000000", "0000000000000111", "0000000000000111"), -- i=28
      ("01", "0000000000000000", "0000000000000111", "1111111111111001"), -- i=29
      ("10", "0000000000000000", "0000000000000111", "0000000000000000"), -- i=30
      ("11", "0000000000000000", "0000000000000111", "0000000000000111"), -- i=31
      ("00", "0000000000000000", "0000000000001000", "0000000000001000"), -- i=32
      ("01", "0000000000000000", "0000000000001000", "1111111111111000"), -- i=33
      ("10", "0000000000000000", "0000000000001000", "0000000000000000"), -- i=34
      ("11", "0000000000000000", "0000000000001000", "0000000000001000"), -- i=35
      ("00", "0000000000000000", "0000000000001001", "0000000000001001"), -- i=36
      ("01", "0000000000000000", "0000000000001001", "1111111111110111"), -- i=37
      ("10", "0000000000000000", "0000000000001001", "0000000000000000"), -- i=38
      ("11", "0000000000000000", "0000000000001001", "0000000000001001"), -- i=39
      ("00", "0000000000000000", "0000000000001010", "0000000000001010"), -- i=40
      ("01", "0000000000000000", "0000000000001010", "1111111111110110"), -- i=41
      ("10", "0000000000000000", "0000000000001010", "0000000000000000"), -- i=42
      ("11", "0000000000000000", "0000000000001010", "0000000000001010"), -- i=43
      ("00", "0000000000000000", "0000000000001011", "0000000000001011"), -- i=44
      ("01", "0000000000000000", "0000000000001011", "1111111111110101"), -- i=45
      ("10", "0000000000000000", "0000000000001011", "0000000000000000"), -- i=46
      ("11", "0000000000000000", "0000000000001011", "0000000000001011"), -- i=47
      ("00", "0000000000000000", "0000000000001100", "0000000000001100"), -- i=48
      ("01", "0000000000000000", "0000000000001100", "1111111111110100"), -- i=49
      ("10", "0000000000000000", "0000000000001100", "0000000000000000"), -- i=50
      ("11", "0000000000000000", "0000000000001100", "0000000000001100"), -- i=51
      ("00", "0000000000000000", "0000000000001101", "0000000000001101"), -- i=52
      ("01", "0000000000000000", "0000000000001101", "1111111111110011"), -- i=53
      ("10", "0000000000000000", "0000000000001101", "0000000000000000"), -- i=54
      ("11", "0000000000000000", "0000000000001101", "0000000000001101"), -- i=55
      ("00", "0000000000000000", "0000000000001110", "0000000000001110"), -- i=56
      ("01", "0000000000000000", "0000000000001110", "1111111111110010"), -- i=57
      ("10", "0000000000000000", "0000000000001110", "0000000000000000"), -- i=58
      ("11", "0000000000000000", "0000000000001110", "0000000000001110"), -- i=59
      ("00", "0000000000000000", "0000000000001111", "0000000000001111"), -- i=60
      ("01", "0000000000000000", "0000000000001111", "1111111111110001"), -- i=61
      ("10", "0000000000000000", "0000000000001111", "0000000000000000"), -- i=62
      ("11", "0000000000000000", "0000000000001111", "0000000000001111"), -- i=63
      ("00", "0000000000000001", "0000000000000000", "0000000000000001"), -- i=64
      ("01", "0000000000000001", "0000000000000000", "0000000000000001"), -- i=65
      ("10", "0000000000000001", "0000000000000000", "0000000000000000"), -- i=66
      ("11", "0000000000000001", "0000000000000000", "0000000000000001"), -- i=67
      ("00", "0000000000000001", "0000000000000001", "0000000000000010"), -- i=68
      ("01", "0000000000000001", "0000000000000001", "0000000000000000"), -- i=69
      ("10", "0000000000000001", "0000000000000001", "0000000000000001"), -- i=70
      ("11", "0000000000000001", "0000000000000001", "0000000000000001"), -- i=71
      ("00", "0000000000000001", "0000000000000010", "0000000000000011"), -- i=72
      ("01", "0000000000000001", "0000000000000010", "1111111111111111"), -- i=73
      ("10", "0000000000000001", "0000000000000010", "0000000000000000"), -- i=74
      ("11", "0000000000000001", "0000000000000010", "0000000000000011"), -- i=75
      ("00", "0000000000000001", "0000000000000011", "0000000000000100"), -- i=76
      ("01", "0000000000000001", "0000000000000011", "1111111111111110"), -- i=77
      ("10", "0000000000000001", "0000000000000011", "0000000000000001"), -- i=78
      ("11", "0000000000000001", "0000000000000011", "0000000000000011"), -- i=79
      ("00", "0000000000000001", "0000000000000100", "0000000000000101"), -- i=80
      ("01", "0000000000000001", "0000000000000100", "1111111111111101"), -- i=81
      ("10", "0000000000000001", "0000000000000100", "0000000000000000"), -- i=82
      ("11", "0000000000000001", "0000000000000100", "0000000000000101"), -- i=83
      ("00", "0000000000000001", "0000000000000101", "0000000000000110"), -- i=84
      ("01", "0000000000000001", "0000000000000101", "1111111111111100"), -- i=85
      ("10", "0000000000000001", "0000000000000101", "0000000000000001"), -- i=86
      ("11", "0000000000000001", "0000000000000101", "0000000000000101"), -- i=87
      ("00", "0000000000000001", "0000000000000110", "0000000000000111"), -- i=88
      ("01", "0000000000000001", "0000000000000110", "1111111111111011"), -- i=89
      ("10", "0000000000000001", "0000000000000110", "0000000000000000"), -- i=90
      ("11", "0000000000000001", "0000000000000110", "0000000000000111"), -- i=91
      ("00", "0000000000000001", "0000000000000111", "0000000000001000"), -- i=92
      ("01", "0000000000000001", "0000000000000111", "1111111111111010"), -- i=93
      ("10", "0000000000000001", "0000000000000111", "0000000000000001"), -- i=94
      ("11", "0000000000000001", "0000000000000111", "0000000000000111"), -- i=95
      ("00", "0000000000000001", "0000000000001000", "0000000000001001"), -- i=96
      ("01", "0000000000000001", "0000000000001000", "1111111111111001"), -- i=97
      ("10", "0000000000000001", "0000000000001000", "0000000000000000"), -- i=98
      ("11", "0000000000000001", "0000000000001000", "0000000000001001"), -- i=99
      ("00", "0000000000000001", "0000000000001001", "0000000000001010"), -- i=100
      ("01", "0000000000000001", "0000000000001001", "1111111111111000"), -- i=101
      ("10", "0000000000000001", "0000000000001001", "0000000000000001"), -- i=102
      ("11", "0000000000000001", "0000000000001001", "0000000000001001"), -- i=103
      ("00", "0000000000000001", "0000000000001010", "0000000000001011"), -- i=104
      ("01", "0000000000000001", "0000000000001010", "1111111111110111"), -- i=105
      ("10", "0000000000000001", "0000000000001010", "0000000000000000"), -- i=106
      ("11", "0000000000000001", "0000000000001010", "0000000000001011"), -- i=107
      ("00", "0000000000000001", "0000000000001011", "0000000000001100"), -- i=108
      ("01", "0000000000000001", "0000000000001011", "1111111111110110"), -- i=109
      ("10", "0000000000000001", "0000000000001011", "0000000000000001"), -- i=110
      ("11", "0000000000000001", "0000000000001011", "0000000000001011"), -- i=111
      ("00", "0000000000000001", "0000000000001100", "0000000000001101"), -- i=112
      ("01", "0000000000000001", "0000000000001100", "1111111111110101"), -- i=113
      ("10", "0000000000000001", "0000000000001100", "0000000000000000"), -- i=114
      ("11", "0000000000000001", "0000000000001100", "0000000000001101"), -- i=115
      ("00", "0000000000000001", "0000000000001101", "0000000000001110"), -- i=116
      ("01", "0000000000000001", "0000000000001101", "1111111111110100"), -- i=117
      ("10", "0000000000000001", "0000000000001101", "0000000000000001"), -- i=118
      ("11", "0000000000000001", "0000000000001101", "0000000000001101"), -- i=119
      ("00", "0000000000000001", "0000000000001110", "0000000000001111"), -- i=120
      ("01", "0000000000000001", "0000000000001110", "1111111111110011"), -- i=121
      ("10", "0000000000000001", "0000000000001110", "0000000000000000"), -- i=122
      ("11", "0000000000000001", "0000000000001110", "0000000000001111"), -- i=123
      ("00", "0000000000000001", "0000000000001111", "0000000000010000"), -- i=124
      ("01", "0000000000000001", "0000000000001111", "1111111111110010"), -- i=125
      ("10", "0000000000000001", "0000000000001111", "0000000000000001"), -- i=126
      ("11", "0000000000000001", "0000000000001111", "0000000000001111"), -- i=127
      ("00", "0000000000000010", "0000000000000000", "0000000000000010"), -- i=128
      ("01", "0000000000000010", "0000000000000000", "0000000000000010"), -- i=129
      ("10", "0000000000000010", "0000000000000000", "0000000000000000"), -- i=130
      ("11", "0000000000000010", "0000000000000000", "0000000000000010"), -- i=131
      ("00", "0000000000000010", "0000000000000001", "0000000000000011"), -- i=132
      ("01", "0000000000000010", "0000000000000001", "0000000000000001"), -- i=133
      ("10", "0000000000000010", "0000000000000001", "0000000000000000"), -- i=134
      ("11", "0000000000000010", "0000000000000001", "0000000000000011"), -- i=135
      ("00", "0000000000000010", "0000000000000010", "0000000000000100"), -- i=136
      ("01", "0000000000000010", "0000000000000010", "0000000000000000"), -- i=137
      ("10", "0000000000000010", "0000000000000010", "0000000000000010"), -- i=138
      ("11", "0000000000000010", "0000000000000010", "0000000000000010"), -- i=139
      ("00", "0000000000000010", "0000000000000011", "0000000000000101"), -- i=140
      ("01", "0000000000000010", "0000000000000011", "1111111111111111"), -- i=141
      ("10", "0000000000000010", "0000000000000011", "0000000000000010"), -- i=142
      ("11", "0000000000000010", "0000000000000011", "0000000000000011"), -- i=143
      ("00", "0000000000000010", "0000000000000100", "0000000000000110"), -- i=144
      ("01", "0000000000000010", "0000000000000100", "1111111111111110"), -- i=145
      ("10", "0000000000000010", "0000000000000100", "0000000000000000"), -- i=146
      ("11", "0000000000000010", "0000000000000100", "0000000000000110"), -- i=147
      ("00", "0000000000000010", "0000000000000101", "0000000000000111"), -- i=148
      ("01", "0000000000000010", "0000000000000101", "1111111111111101"), -- i=149
      ("10", "0000000000000010", "0000000000000101", "0000000000000000"), -- i=150
      ("11", "0000000000000010", "0000000000000101", "0000000000000111"), -- i=151
      ("00", "0000000000000010", "0000000000000110", "0000000000001000"), -- i=152
      ("01", "0000000000000010", "0000000000000110", "1111111111111100"), -- i=153
      ("10", "0000000000000010", "0000000000000110", "0000000000000010"), -- i=154
      ("11", "0000000000000010", "0000000000000110", "0000000000000110"), -- i=155
      ("00", "0000000000000010", "0000000000000111", "0000000000001001"), -- i=156
      ("01", "0000000000000010", "0000000000000111", "1111111111111011"), -- i=157
      ("10", "0000000000000010", "0000000000000111", "0000000000000010"), -- i=158
      ("11", "0000000000000010", "0000000000000111", "0000000000000111"), -- i=159
      ("00", "0000000000000010", "0000000000001000", "0000000000001010"), -- i=160
      ("01", "0000000000000010", "0000000000001000", "1111111111111010"), -- i=161
      ("10", "0000000000000010", "0000000000001000", "0000000000000000"), -- i=162
      ("11", "0000000000000010", "0000000000001000", "0000000000001010"), -- i=163
      ("00", "0000000000000010", "0000000000001001", "0000000000001011"), -- i=164
      ("01", "0000000000000010", "0000000000001001", "1111111111111001"), -- i=165
      ("10", "0000000000000010", "0000000000001001", "0000000000000000"), -- i=166
      ("11", "0000000000000010", "0000000000001001", "0000000000001011"), -- i=167
      ("00", "0000000000000010", "0000000000001010", "0000000000001100"), -- i=168
      ("01", "0000000000000010", "0000000000001010", "1111111111111000"), -- i=169
      ("10", "0000000000000010", "0000000000001010", "0000000000000010"), -- i=170
      ("11", "0000000000000010", "0000000000001010", "0000000000001010"), -- i=171
      ("00", "0000000000000010", "0000000000001011", "0000000000001101"), -- i=172
      ("01", "0000000000000010", "0000000000001011", "1111111111110111"), -- i=173
      ("10", "0000000000000010", "0000000000001011", "0000000000000010"), -- i=174
      ("11", "0000000000000010", "0000000000001011", "0000000000001011"), -- i=175
      ("00", "0000000000000010", "0000000000001100", "0000000000001110"), -- i=176
      ("01", "0000000000000010", "0000000000001100", "1111111111110110"), -- i=177
      ("10", "0000000000000010", "0000000000001100", "0000000000000000"), -- i=178
      ("11", "0000000000000010", "0000000000001100", "0000000000001110"), -- i=179
      ("00", "0000000000000010", "0000000000001101", "0000000000001111"), -- i=180
      ("01", "0000000000000010", "0000000000001101", "1111111111110101"), -- i=181
      ("10", "0000000000000010", "0000000000001101", "0000000000000000"), -- i=182
      ("11", "0000000000000010", "0000000000001101", "0000000000001111"), -- i=183
      ("00", "0000000000000010", "0000000000001110", "0000000000010000"), -- i=184
      ("01", "0000000000000010", "0000000000001110", "1111111111110100"), -- i=185
      ("10", "0000000000000010", "0000000000001110", "0000000000000010"), -- i=186
      ("11", "0000000000000010", "0000000000001110", "0000000000001110"), -- i=187
      ("00", "0000000000000010", "0000000000001111", "0000000000010001"), -- i=188
      ("01", "0000000000000010", "0000000000001111", "1111111111110011"), -- i=189
      ("10", "0000000000000010", "0000000000001111", "0000000000000010"), -- i=190
      ("11", "0000000000000010", "0000000000001111", "0000000000001111"), -- i=191
      ("00", "0000000000000011", "0000000000000000", "0000000000000011"), -- i=192
      ("01", "0000000000000011", "0000000000000000", "0000000000000011"), -- i=193
      ("10", "0000000000000011", "0000000000000000", "0000000000000000"), -- i=194
      ("11", "0000000000000011", "0000000000000000", "0000000000000011"), -- i=195
      ("00", "0000000000000011", "0000000000000001", "0000000000000100"), -- i=196
      ("01", "0000000000000011", "0000000000000001", "0000000000000010"), -- i=197
      ("10", "0000000000000011", "0000000000000001", "0000000000000001"), -- i=198
      ("11", "0000000000000011", "0000000000000001", "0000000000000011"), -- i=199
      ("00", "0000000000000011", "0000000000000010", "0000000000000101"), -- i=200
      ("01", "0000000000000011", "0000000000000010", "0000000000000001"), -- i=201
      ("10", "0000000000000011", "0000000000000010", "0000000000000010"), -- i=202
      ("11", "0000000000000011", "0000000000000010", "0000000000000011"), -- i=203
      ("00", "0000000000000011", "0000000000000011", "0000000000000110"), -- i=204
      ("01", "0000000000000011", "0000000000000011", "0000000000000000"), -- i=205
      ("10", "0000000000000011", "0000000000000011", "0000000000000011"), -- i=206
      ("11", "0000000000000011", "0000000000000011", "0000000000000011"), -- i=207
      ("00", "0000000000000011", "0000000000000100", "0000000000000111"), -- i=208
      ("01", "0000000000000011", "0000000000000100", "1111111111111111"), -- i=209
      ("10", "0000000000000011", "0000000000000100", "0000000000000000"), -- i=210
      ("11", "0000000000000011", "0000000000000100", "0000000000000111"), -- i=211
      ("00", "0000000000000011", "0000000000000101", "0000000000001000"), -- i=212
      ("01", "0000000000000011", "0000000000000101", "1111111111111110"), -- i=213
      ("10", "0000000000000011", "0000000000000101", "0000000000000001"), -- i=214
      ("11", "0000000000000011", "0000000000000101", "0000000000000111"), -- i=215
      ("00", "0000000000000011", "0000000000000110", "0000000000001001"), -- i=216
      ("01", "0000000000000011", "0000000000000110", "1111111111111101"), -- i=217
      ("10", "0000000000000011", "0000000000000110", "0000000000000010"), -- i=218
      ("11", "0000000000000011", "0000000000000110", "0000000000000111"), -- i=219
      ("00", "0000000000000011", "0000000000000111", "0000000000001010"), -- i=220
      ("01", "0000000000000011", "0000000000000111", "1111111111111100"), -- i=221
      ("10", "0000000000000011", "0000000000000111", "0000000000000011"), -- i=222
      ("11", "0000000000000011", "0000000000000111", "0000000000000111"), -- i=223
      ("00", "0000000000000011", "0000000000001000", "0000000000001011"), -- i=224
      ("01", "0000000000000011", "0000000000001000", "1111111111111011"), -- i=225
      ("10", "0000000000000011", "0000000000001000", "0000000000000000"), -- i=226
      ("11", "0000000000000011", "0000000000001000", "0000000000001011"), -- i=227
      ("00", "0000000000000011", "0000000000001001", "0000000000001100"), -- i=228
      ("01", "0000000000000011", "0000000000001001", "1111111111111010"), -- i=229
      ("10", "0000000000000011", "0000000000001001", "0000000000000001"), -- i=230
      ("11", "0000000000000011", "0000000000001001", "0000000000001011"), -- i=231
      ("00", "0000000000000011", "0000000000001010", "0000000000001101"), -- i=232
      ("01", "0000000000000011", "0000000000001010", "1111111111111001"), -- i=233
      ("10", "0000000000000011", "0000000000001010", "0000000000000010"), -- i=234
      ("11", "0000000000000011", "0000000000001010", "0000000000001011"), -- i=235
      ("00", "0000000000000011", "0000000000001011", "0000000000001110"), -- i=236
      ("01", "0000000000000011", "0000000000001011", "1111111111111000"), -- i=237
      ("10", "0000000000000011", "0000000000001011", "0000000000000011"), -- i=238
      ("11", "0000000000000011", "0000000000001011", "0000000000001011"), -- i=239
      ("00", "0000000000000011", "0000000000001100", "0000000000001111"), -- i=240
      ("01", "0000000000000011", "0000000000001100", "1111111111110111"), -- i=241
      ("10", "0000000000000011", "0000000000001100", "0000000000000000"), -- i=242
      ("11", "0000000000000011", "0000000000001100", "0000000000001111"), -- i=243
      ("00", "0000000000000011", "0000000000001101", "0000000000010000"), -- i=244
      ("01", "0000000000000011", "0000000000001101", "1111111111110110"), -- i=245
      ("10", "0000000000000011", "0000000000001101", "0000000000000001"), -- i=246
      ("11", "0000000000000011", "0000000000001101", "0000000000001111"), -- i=247
      ("00", "0000000000000011", "0000000000001110", "0000000000010001"), -- i=248
      ("01", "0000000000000011", "0000000000001110", "1111111111110101"), -- i=249
      ("10", "0000000000000011", "0000000000001110", "0000000000000010"), -- i=250
      ("11", "0000000000000011", "0000000000001110", "0000000000001111"), -- i=251
      ("00", "0000000000000011", "0000000000001111", "0000000000010010"), -- i=252
      ("01", "0000000000000011", "0000000000001111", "1111111111110100"), -- i=253
      ("10", "0000000000000011", "0000000000001111", "0000000000000011"), -- i=254
      ("11", "0000000000000011", "0000000000001111", "0000000000001111"), -- i=255
      ("00", "0000000000000100", "0000000000000000", "0000000000000100"), -- i=256
      ("01", "0000000000000100", "0000000000000000", "0000000000000100"), -- i=257
      ("10", "0000000000000100", "0000000000000000", "0000000000000000"), -- i=258
      ("11", "0000000000000100", "0000000000000000", "0000000000000100"), -- i=259
      ("00", "0000000000000100", "0000000000000001", "0000000000000101"), -- i=260
      ("01", "0000000000000100", "0000000000000001", "0000000000000011"), -- i=261
      ("10", "0000000000000100", "0000000000000001", "0000000000000000"), -- i=262
      ("11", "0000000000000100", "0000000000000001", "0000000000000101"), -- i=263
      ("00", "0000000000000100", "0000000000000010", "0000000000000110"), -- i=264
      ("01", "0000000000000100", "0000000000000010", "0000000000000010"), -- i=265
      ("10", "0000000000000100", "0000000000000010", "0000000000000000"), -- i=266
      ("11", "0000000000000100", "0000000000000010", "0000000000000110"), -- i=267
      ("00", "0000000000000100", "0000000000000011", "0000000000000111"), -- i=268
      ("01", "0000000000000100", "0000000000000011", "0000000000000001"), -- i=269
      ("10", "0000000000000100", "0000000000000011", "0000000000000000"), -- i=270
      ("11", "0000000000000100", "0000000000000011", "0000000000000111"), -- i=271
      ("00", "0000000000000100", "0000000000000100", "0000000000001000"), -- i=272
      ("01", "0000000000000100", "0000000000000100", "0000000000000000"), -- i=273
      ("10", "0000000000000100", "0000000000000100", "0000000000000100"), -- i=274
      ("11", "0000000000000100", "0000000000000100", "0000000000000100"), -- i=275
      ("00", "0000000000000100", "0000000000000101", "0000000000001001"), -- i=276
      ("01", "0000000000000100", "0000000000000101", "1111111111111111"), -- i=277
      ("10", "0000000000000100", "0000000000000101", "0000000000000100"), -- i=278
      ("11", "0000000000000100", "0000000000000101", "0000000000000101"), -- i=279
      ("00", "0000000000000100", "0000000000000110", "0000000000001010"), -- i=280
      ("01", "0000000000000100", "0000000000000110", "1111111111111110"), -- i=281
      ("10", "0000000000000100", "0000000000000110", "0000000000000100"), -- i=282
      ("11", "0000000000000100", "0000000000000110", "0000000000000110"), -- i=283
      ("00", "0000000000000100", "0000000000000111", "0000000000001011"), -- i=284
      ("01", "0000000000000100", "0000000000000111", "1111111111111101"), -- i=285
      ("10", "0000000000000100", "0000000000000111", "0000000000000100"), -- i=286
      ("11", "0000000000000100", "0000000000000111", "0000000000000111"), -- i=287
      ("00", "0000000000000100", "0000000000001000", "0000000000001100"), -- i=288
      ("01", "0000000000000100", "0000000000001000", "1111111111111100"), -- i=289
      ("10", "0000000000000100", "0000000000001000", "0000000000000000"), -- i=290
      ("11", "0000000000000100", "0000000000001000", "0000000000001100"), -- i=291
      ("00", "0000000000000100", "0000000000001001", "0000000000001101"), -- i=292
      ("01", "0000000000000100", "0000000000001001", "1111111111111011"), -- i=293
      ("10", "0000000000000100", "0000000000001001", "0000000000000000"), -- i=294
      ("11", "0000000000000100", "0000000000001001", "0000000000001101"), -- i=295
      ("00", "0000000000000100", "0000000000001010", "0000000000001110"), -- i=296
      ("01", "0000000000000100", "0000000000001010", "1111111111111010"), -- i=297
      ("10", "0000000000000100", "0000000000001010", "0000000000000000"), -- i=298
      ("11", "0000000000000100", "0000000000001010", "0000000000001110"), -- i=299
      ("00", "0000000000000100", "0000000000001011", "0000000000001111"), -- i=300
      ("01", "0000000000000100", "0000000000001011", "1111111111111001"), -- i=301
      ("10", "0000000000000100", "0000000000001011", "0000000000000000"), -- i=302
      ("11", "0000000000000100", "0000000000001011", "0000000000001111"), -- i=303
      ("00", "0000000000000100", "0000000000001100", "0000000000010000"), -- i=304
      ("01", "0000000000000100", "0000000000001100", "1111111111111000"), -- i=305
      ("10", "0000000000000100", "0000000000001100", "0000000000000100"), -- i=306
      ("11", "0000000000000100", "0000000000001100", "0000000000001100"), -- i=307
      ("00", "0000000000000100", "0000000000001101", "0000000000010001"), -- i=308
      ("01", "0000000000000100", "0000000000001101", "1111111111110111"), -- i=309
      ("10", "0000000000000100", "0000000000001101", "0000000000000100"), -- i=310
      ("11", "0000000000000100", "0000000000001101", "0000000000001101"), -- i=311
      ("00", "0000000000000100", "0000000000001110", "0000000000010010"), -- i=312
      ("01", "0000000000000100", "0000000000001110", "1111111111110110"), -- i=313
      ("10", "0000000000000100", "0000000000001110", "0000000000000100"), -- i=314
      ("11", "0000000000000100", "0000000000001110", "0000000000001110"), -- i=315
      ("00", "0000000000000100", "0000000000001111", "0000000000010011"), -- i=316
      ("01", "0000000000000100", "0000000000001111", "1111111111110101"), -- i=317
      ("10", "0000000000000100", "0000000000001111", "0000000000000100"), -- i=318
      ("11", "0000000000000100", "0000000000001111", "0000000000001111"), -- i=319
      ("00", "0000000000000101", "0000000000000000", "0000000000000101"), -- i=320
      ("01", "0000000000000101", "0000000000000000", "0000000000000101"), -- i=321
      ("10", "0000000000000101", "0000000000000000", "0000000000000000"), -- i=322
      ("11", "0000000000000101", "0000000000000000", "0000000000000101"), -- i=323
      ("00", "0000000000000101", "0000000000000001", "0000000000000110"), -- i=324
      ("01", "0000000000000101", "0000000000000001", "0000000000000100"), -- i=325
      ("10", "0000000000000101", "0000000000000001", "0000000000000001"), -- i=326
      ("11", "0000000000000101", "0000000000000001", "0000000000000101"), -- i=327
      ("00", "0000000000000101", "0000000000000010", "0000000000000111"), -- i=328
      ("01", "0000000000000101", "0000000000000010", "0000000000000011"), -- i=329
      ("10", "0000000000000101", "0000000000000010", "0000000000000000"), -- i=330
      ("11", "0000000000000101", "0000000000000010", "0000000000000111"), -- i=331
      ("00", "0000000000000101", "0000000000000011", "0000000000001000"), -- i=332
      ("01", "0000000000000101", "0000000000000011", "0000000000000010"), -- i=333
      ("10", "0000000000000101", "0000000000000011", "0000000000000001"), -- i=334
      ("11", "0000000000000101", "0000000000000011", "0000000000000111"), -- i=335
      ("00", "0000000000000101", "0000000000000100", "0000000000001001"), -- i=336
      ("01", "0000000000000101", "0000000000000100", "0000000000000001"), -- i=337
      ("10", "0000000000000101", "0000000000000100", "0000000000000100"), -- i=338
      ("11", "0000000000000101", "0000000000000100", "0000000000000101"), -- i=339
      ("00", "0000000000000101", "0000000000000101", "0000000000001010"), -- i=340
      ("01", "0000000000000101", "0000000000000101", "0000000000000000"), -- i=341
      ("10", "0000000000000101", "0000000000000101", "0000000000000101"), -- i=342
      ("11", "0000000000000101", "0000000000000101", "0000000000000101"), -- i=343
      ("00", "0000000000000101", "0000000000000110", "0000000000001011"), -- i=344
      ("01", "0000000000000101", "0000000000000110", "1111111111111111"), -- i=345
      ("10", "0000000000000101", "0000000000000110", "0000000000000100"), -- i=346
      ("11", "0000000000000101", "0000000000000110", "0000000000000111"), -- i=347
      ("00", "0000000000000101", "0000000000000111", "0000000000001100"), -- i=348
      ("01", "0000000000000101", "0000000000000111", "1111111111111110"), -- i=349
      ("10", "0000000000000101", "0000000000000111", "0000000000000101"), -- i=350
      ("11", "0000000000000101", "0000000000000111", "0000000000000111"), -- i=351
      ("00", "0000000000000101", "0000000000001000", "0000000000001101"), -- i=352
      ("01", "0000000000000101", "0000000000001000", "1111111111111101"), -- i=353
      ("10", "0000000000000101", "0000000000001000", "0000000000000000"), -- i=354
      ("11", "0000000000000101", "0000000000001000", "0000000000001101"), -- i=355
      ("00", "0000000000000101", "0000000000001001", "0000000000001110"), -- i=356
      ("01", "0000000000000101", "0000000000001001", "1111111111111100"), -- i=357
      ("10", "0000000000000101", "0000000000001001", "0000000000000001"), -- i=358
      ("11", "0000000000000101", "0000000000001001", "0000000000001101"), -- i=359
      ("00", "0000000000000101", "0000000000001010", "0000000000001111"), -- i=360
      ("01", "0000000000000101", "0000000000001010", "1111111111111011"), -- i=361
      ("10", "0000000000000101", "0000000000001010", "0000000000000000"), -- i=362
      ("11", "0000000000000101", "0000000000001010", "0000000000001111"), -- i=363
      ("00", "0000000000000101", "0000000000001011", "0000000000010000"), -- i=364
      ("01", "0000000000000101", "0000000000001011", "1111111111111010"), -- i=365
      ("10", "0000000000000101", "0000000000001011", "0000000000000001"), -- i=366
      ("11", "0000000000000101", "0000000000001011", "0000000000001111"), -- i=367
      ("00", "0000000000000101", "0000000000001100", "0000000000010001"), -- i=368
      ("01", "0000000000000101", "0000000000001100", "1111111111111001"), -- i=369
      ("10", "0000000000000101", "0000000000001100", "0000000000000100"), -- i=370
      ("11", "0000000000000101", "0000000000001100", "0000000000001101"), -- i=371
      ("00", "0000000000000101", "0000000000001101", "0000000000010010"), -- i=372
      ("01", "0000000000000101", "0000000000001101", "1111111111111000"), -- i=373
      ("10", "0000000000000101", "0000000000001101", "0000000000000101"), -- i=374
      ("11", "0000000000000101", "0000000000001101", "0000000000001101"), -- i=375
      ("00", "0000000000000101", "0000000000001110", "0000000000010011"), -- i=376
      ("01", "0000000000000101", "0000000000001110", "1111111111110111"), -- i=377
      ("10", "0000000000000101", "0000000000001110", "0000000000000100"), -- i=378
      ("11", "0000000000000101", "0000000000001110", "0000000000001111"), -- i=379
      ("00", "0000000000000101", "0000000000001111", "0000000000010100"), -- i=380
      ("01", "0000000000000101", "0000000000001111", "1111111111110110"), -- i=381
      ("10", "0000000000000101", "0000000000001111", "0000000000000101"), -- i=382
      ("11", "0000000000000101", "0000000000001111", "0000000000001111"), -- i=383
      ("00", "0000000000000110", "0000000000000000", "0000000000000110"), -- i=384
      ("01", "0000000000000110", "0000000000000000", "0000000000000110"), -- i=385
      ("10", "0000000000000110", "0000000000000000", "0000000000000000"), -- i=386
      ("11", "0000000000000110", "0000000000000000", "0000000000000110"), -- i=387
      ("00", "0000000000000110", "0000000000000001", "0000000000000111"), -- i=388
      ("01", "0000000000000110", "0000000000000001", "0000000000000101"), -- i=389
      ("10", "0000000000000110", "0000000000000001", "0000000000000000"), -- i=390
      ("11", "0000000000000110", "0000000000000001", "0000000000000111"), -- i=391
      ("00", "0000000000000110", "0000000000000010", "0000000000001000"), -- i=392
      ("01", "0000000000000110", "0000000000000010", "0000000000000100"), -- i=393
      ("10", "0000000000000110", "0000000000000010", "0000000000000010"), -- i=394
      ("11", "0000000000000110", "0000000000000010", "0000000000000110"), -- i=395
      ("00", "0000000000000110", "0000000000000011", "0000000000001001"), -- i=396
      ("01", "0000000000000110", "0000000000000011", "0000000000000011"), -- i=397
      ("10", "0000000000000110", "0000000000000011", "0000000000000010"), -- i=398
      ("11", "0000000000000110", "0000000000000011", "0000000000000111"), -- i=399
      ("00", "0000000000000110", "0000000000000100", "0000000000001010"), -- i=400
      ("01", "0000000000000110", "0000000000000100", "0000000000000010"), -- i=401
      ("10", "0000000000000110", "0000000000000100", "0000000000000100"), -- i=402
      ("11", "0000000000000110", "0000000000000100", "0000000000000110"), -- i=403
      ("00", "0000000000000110", "0000000000000101", "0000000000001011"), -- i=404
      ("01", "0000000000000110", "0000000000000101", "0000000000000001"), -- i=405
      ("10", "0000000000000110", "0000000000000101", "0000000000000100"), -- i=406
      ("11", "0000000000000110", "0000000000000101", "0000000000000111"), -- i=407
      ("00", "0000000000000110", "0000000000000110", "0000000000001100"), -- i=408
      ("01", "0000000000000110", "0000000000000110", "0000000000000000"), -- i=409
      ("10", "0000000000000110", "0000000000000110", "0000000000000110"), -- i=410
      ("11", "0000000000000110", "0000000000000110", "0000000000000110"), -- i=411
      ("00", "0000000000000110", "0000000000000111", "0000000000001101"), -- i=412
      ("01", "0000000000000110", "0000000000000111", "1111111111111111"), -- i=413
      ("10", "0000000000000110", "0000000000000111", "0000000000000110"), -- i=414
      ("11", "0000000000000110", "0000000000000111", "0000000000000111"), -- i=415
      ("00", "0000000000000110", "0000000000001000", "0000000000001110"), -- i=416
      ("01", "0000000000000110", "0000000000001000", "1111111111111110"), -- i=417
      ("10", "0000000000000110", "0000000000001000", "0000000000000000"), -- i=418
      ("11", "0000000000000110", "0000000000001000", "0000000000001110"), -- i=419
      ("00", "0000000000000110", "0000000000001001", "0000000000001111"), -- i=420
      ("01", "0000000000000110", "0000000000001001", "1111111111111101"), -- i=421
      ("10", "0000000000000110", "0000000000001001", "0000000000000000"), -- i=422
      ("11", "0000000000000110", "0000000000001001", "0000000000001111"), -- i=423
      ("00", "0000000000000110", "0000000000001010", "0000000000010000"), -- i=424
      ("01", "0000000000000110", "0000000000001010", "1111111111111100"), -- i=425
      ("10", "0000000000000110", "0000000000001010", "0000000000000010"), -- i=426
      ("11", "0000000000000110", "0000000000001010", "0000000000001110"), -- i=427
      ("00", "0000000000000110", "0000000000001011", "0000000000010001"), -- i=428
      ("01", "0000000000000110", "0000000000001011", "1111111111111011"), -- i=429
      ("10", "0000000000000110", "0000000000001011", "0000000000000010"), -- i=430
      ("11", "0000000000000110", "0000000000001011", "0000000000001111"), -- i=431
      ("00", "0000000000000110", "0000000000001100", "0000000000010010"), -- i=432
      ("01", "0000000000000110", "0000000000001100", "1111111111111010"), -- i=433
      ("10", "0000000000000110", "0000000000001100", "0000000000000100"), -- i=434
      ("11", "0000000000000110", "0000000000001100", "0000000000001110"), -- i=435
      ("00", "0000000000000110", "0000000000001101", "0000000000010011"), -- i=436
      ("01", "0000000000000110", "0000000000001101", "1111111111111001"), -- i=437
      ("10", "0000000000000110", "0000000000001101", "0000000000000100"), -- i=438
      ("11", "0000000000000110", "0000000000001101", "0000000000001111"), -- i=439
      ("00", "0000000000000110", "0000000000001110", "0000000000010100"), -- i=440
      ("01", "0000000000000110", "0000000000001110", "1111111111111000"), -- i=441
      ("10", "0000000000000110", "0000000000001110", "0000000000000110"), -- i=442
      ("11", "0000000000000110", "0000000000001110", "0000000000001110"), -- i=443
      ("00", "0000000000000110", "0000000000001111", "0000000000010101"), -- i=444
      ("01", "0000000000000110", "0000000000001111", "1111111111110111"), -- i=445
      ("10", "0000000000000110", "0000000000001111", "0000000000000110"), -- i=446
      ("11", "0000000000000110", "0000000000001111", "0000000000001111"), -- i=447
      ("00", "0000000000000111", "0000000000000000", "0000000000000111"), -- i=448
      ("01", "0000000000000111", "0000000000000000", "0000000000000111"), -- i=449
      ("10", "0000000000000111", "0000000000000000", "0000000000000000"), -- i=450
      ("11", "0000000000000111", "0000000000000000", "0000000000000111"), -- i=451
      ("00", "0000000000000111", "0000000000000001", "0000000000001000"), -- i=452
      ("01", "0000000000000111", "0000000000000001", "0000000000000110"), -- i=453
      ("10", "0000000000000111", "0000000000000001", "0000000000000001"), -- i=454
      ("11", "0000000000000111", "0000000000000001", "0000000000000111"), -- i=455
      ("00", "0000000000000111", "0000000000000010", "0000000000001001"), -- i=456
      ("01", "0000000000000111", "0000000000000010", "0000000000000101"), -- i=457
      ("10", "0000000000000111", "0000000000000010", "0000000000000010"), -- i=458
      ("11", "0000000000000111", "0000000000000010", "0000000000000111"), -- i=459
      ("00", "0000000000000111", "0000000000000011", "0000000000001010"), -- i=460
      ("01", "0000000000000111", "0000000000000011", "0000000000000100"), -- i=461
      ("10", "0000000000000111", "0000000000000011", "0000000000000011"), -- i=462
      ("11", "0000000000000111", "0000000000000011", "0000000000000111"), -- i=463
      ("00", "0000000000000111", "0000000000000100", "0000000000001011"), -- i=464
      ("01", "0000000000000111", "0000000000000100", "0000000000000011"), -- i=465
      ("10", "0000000000000111", "0000000000000100", "0000000000000100"), -- i=466
      ("11", "0000000000000111", "0000000000000100", "0000000000000111"), -- i=467
      ("00", "0000000000000111", "0000000000000101", "0000000000001100"), -- i=468
      ("01", "0000000000000111", "0000000000000101", "0000000000000010"), -- i=469
      ("10", "0000000000000111", "0000000000000101", "0000000000000101"), -- i=470
      ("11", "0000000000000111", "0000000000000101", "0000000000000111"), -- i=471
      ("00", "0000000000000111", "0000000000000110", "0000000000001101"), -- i=472
      ("01", "0000000000000111", "0000000000000110", "0000000000000001"), -- i=473
      ("10", "0000000000000111", "0000000000000110", "0000000000000110"), -- i=474
      ("11", "0000000000000111", "0000000000000110", "0000000000000111"), -- i=475
      ("00", "0000000000000111", "0000000000000111", "0000000000001110"), -- i=476
      ("01", "0000000000000111", "0000000000000111", "0000000000000000"), -- i=477
      ("10", "0000000000000111", "0000000000000111", "0000000000000111"), -- i=478
      ("11", "0000000000000111", "0000000000000111", "0000000000000111"), -- i=479
      ("00", "0000000000000111", "0000000000001000", "0000000000001111"), -- i=480
      ("01", "0000000000000111", "0000000000001000", "1111111111111111"), -- i=481
      ("10", "0000000000000111", "0000000000001000", "0000000000000000"), -- i=482
      ("11", "0000000000000111", "0000000000001000", "0000000000001111"), -- i=483
      ("00", "0000000000000111", "0000000000001001", "0000000000010000"), -- i=484
      ("01", "0000000000000111", "0000000000001001", "1111111111111110"), -- i=485
      ("10", "0000000000000111", "0000000000001001", "0000000000000001"), -- i=486
      ("11", "0000000000000111", "0000000000001001", "0000000000001111"), -- i=487
      ("00", "0000000000000111", "0000000000001010", "0000000000010001"), -- i=488
      ("01", "0000000000000111", "0000000000001010", "1111111111111101"), -- i=489
      ("10", "0000000000000111", "0000000000001010", "0000000000000010"), -- i=490
      ("11", "0000000000000111", "0000000000001010", "0000000000001111"), -- i=491
      ("00", "0000000000000111", "0000000000001011", "0000000000010010"), -- i=492
      ("01", "0000000000000111", "0000000000001011", "1111111111111100"), -- i=493
      ("10", "0000000000000111", "0000000000001011", "0000000000000011"), -- i=494
      ("11", "0000000000000111", "0000000000001011", "0000000000001111"), -- i=495
      ("00", "0000000000000111", "0000000000001100", "0000000000010011"), -- i=496
      ("01", "0000000000000111", "0000000000001100", "1111111111111011"), -- i=497
      ("10", "0000000000000111", "0000000000001100", "0000000000000100"), -- i=498
      ("11", "0000000000000111", "0000000000001100", "0000000000001111"), -- i=499
      ("00", "0000000000000111", "0000000000001101", "0000000000010100"), -- i=500
      ("01", "0000000000000111", "0000000000001101", "1111111111111010"), -- i=501
      ("10", "0000000000000111", "0000000000001101", "0000000000000101"), -- i=502
      ("11", "0000000000000111", "0000000000001101", "0000000000001111"), -- i=503
      ("00", "0000000000000111", "0000000000001110", "0000000000010101"), -- i=504
      ("01", "0000000000000111", "0000000000001110", "1111111111111001"), -- i=505
      ("10", "0000000000000111", "0000000000001110", "0000000000000110"), -- i=506
      ("11", "0000000000000111", "0000000000001110", "0000000000001111"), -- i=507
      ("00", "0000000000000111", "0000000000001111", "0000000000010110"), -- i=508
      ("01", "0000000000000111", "0000000000001111", "1111111111111000"), -- i=509
      ("10", "0000000000000111", "0000000000001111", "0000000000000111"), -- i=510
      ("11", "0000000000000111", "0000000000001111", "0000000000001111"), -- i=511
      ("00", "0000000000001000", "0000000000000000", "0000000000001000"), -- i=512
      ("01", "0000000000001000", "0000000000000000", "0000000000001000"), -- i=513
      ("10", "0000000000001000", "0000000000000000", "0000000000000000"), -- i=514
      ("11", "0000000000001000", "0000000000000000", "0000000000001000"), -- i=515
      ("00", "0000000000001000", "0000000000000001", "0000000000001001"), -- i=516
      ("01", "0000000000001000", "0000000000000001", "0000000000000111"), -- i=517
      ("10", "0000000000001000", "0000000000000001", "0000000000000000"), -- i=518
      ("11", "0000000000001000", "0000000000000001", "0000000000001001"), -- i=519
      ("00", "0000000000001000", "0000000000000010", "0000000000001010"), -- i=520
      ("01", "0000000000001000", "0000000000000010", "0000000000000110"), -- i=521
      ("10", "0000000000001000", "0000000000000010", "0000000000000000"), -- i=522
      ("11", "0000000000001000", "0000000000000010", "0000000000001010"), -- i=523
      ("00", "0000000000001000", "0000000000000011", "0000000000001011"), -- i=524
      ("01", "0000000000001000", "0000000000000011", "0000000000000101"), -- i=525
      ("10", "0000000000001000", "0000000000000011", "0000000000000000"), -- i=526
      ("11", "0000000000001000", "0000000000000011", "0000000000001011"), -- i=527
      ("00", "0000000000001000", "0000000000000100", "0000000000001100"), -- i=528
      ("01", "0000000000001000", "0000000000000100", "0000000000000100"), -- i=529
      ("10", "0000000000001000", "0000000000000100", "0000000000000000"), -- i=530
      ("11", "0000000000001000", "0000000000000100", "0000000000001100"), -- i=531
      ("00", "0000000000001000", "0000000000000101", "0000000000001101"), -- i=532
      ("01", "0000000000001000", "0000000000000101", "0000000000000011"), -- i=533
      ("10", "0000000000001000", "0000000000000101", "0000000000000000"), -- i=534
      ("11", "0000000000001000", "0000000000000101", "0000000000001101"), -- i=535
      ("00", "0000000000001000", "0000000000000110", "0000000000001110"), -- i=536
      ("01", "0000000000001000", "0000000000000110", "0000000000000010"), -- i=537
      ("10", "0000000000001000", "0000000000000110", "0000000000000000"), -- i=538
      ("11", "0000000000001000", "0000000000000110", "0000000000001110"), -- i=539
      ("00", "0000000000001000", "0000000000000111", "0000000000001111"), -- i=540
      ("01", "0000000000001000", "0000000000000111", "0000000000000001"), -- i=541
      ("10", "0000000000001000", "0000000000000111", "0000000000000000"), -- i=542
      ("11", "0000000000001000", "0000000000000111", "0000000000001111"), -- i=543
      ("00", "0000000000001000", "0000000000001000", "0000000000010000"), -- i=544
      ("01", "0000000000001000", "0000000000001000", "0000000000000000"), -- i=545
      ("10", "0000000000001000", "0000000000001000", "0000000000001000"), -- i=546
      ("11", "0000000000001000", "0000000000001000", "0000000000001000"), -- i=547
      ("00", "0000000000001000", "0000000000001001", "0000000000010001"), -- i=548
      ("01", "0000000000001000", "0000000000001001", "1111111111111111"), -- i=549
      ("10", "0000000000001000", "0000000000001001", "0000000000001000"), -- i=550
      ("11", "0000000000001000", "0000000000001001", "0000000000001001"), -- i=551
      ("00", "0000000000001000", "0000000000001010", "0000000000010010"), -- i=552
      ("01", "0000000000001000", "0000000000001010", "1111111111111110"), -- i=553
      ("10", "0000000000001000", "0000000000001010", "0000000000001000"), -- i=554
      ("11", "0000000000001000", "0000000000001010", "0000000000001010"), -- i=555
      ("00", "0000000000001000", "0000000000001011", "0000000000010011"), -- i=556
      ("01", "0000000000001000", "0000000000001011", "1111111111111101"), -- i=557
      ("10", "0000000000001000", "0000000000001011", "0000000000001000"), -- i=558
      ("11", "0000000000001000", "0000000000001011", "0000000000001011"), -- i=559
      ("00", "0000000000001000", "0000000000001100", "0000000000010100"), -- i=560
      ("01", "0000000000001000", "0000000000001100", "1111111111111100"), -- i=561
      ("10", "0000000000001000", "0000000000001100", "0000000000001000"), -- i=562
      ("11", "0000000000001000", "0000000000001100", "0000000000001100"), -- i=563
      ("00", "0000000000001000", "0000000000001101", "0000000000010101"), -- i=564
      ("01", "0000000000001000", "0000000000001101", "1111111111111011"), -- i=565
      ("10", "0000000000001000", "0000000000001101", "0000000000001000"), -- i=566
      ("11", "0000000000001000", "0000000000001101", "0000000000001101"), -- i=567
      ("00", "0000000000001000", "0000000000001110", "0000000000010110"), -- i=568
      ("01", "0000000000001000", "0000000000001110", "1111111111111010"), -- i=569
      ("10", "0000000000001000", "0000000000001110", "0000000000001000"), -- i=570
      ("11", "0000000000001000", "0000000000001110", "0000000000001110"), -- i=571
      ("00", "0000000000001000", "0000000000001111", "0000000000010111"), -- i=572
      ("01", "0000000000001000", "0000000000001111", "1111111111111001"), -- i=573
      ("10", "0000000000001000", "0000000000001111", "0000000000001000"), -- i=574
      ("11", "0000000000001000", "0000000000001111", "0000000000001111"), -- i=575
      ("00", "0000000000001001", "0000000000000000", "0000000000001001"), -- i=576
      ("01", "0000000000001001", "0000000000000000", "0000000000001001"), -- i=577
      ("10", "0000000000001001", "0000000000000000", "0000000000000000"), -- i=578
      ("11", "0000000000001001", "0000000000000000", "0000000000001001"), -- i=579
      ("00", "0000000000001001", "0000000000000001", "0000000000001010"), -- i=580
      ("01", "0000000000001001", "0000000000000001", "0000000000001000"), -- i=581
      ("10", "0000000000001001", "0000000000000001", "0000000000000001"), -- i=582
      ("11", "0000000000001001", "0000000000000001", "0000000000001001"), -- i=583
      ("00", "0000000000001001", "0000000000000010", "0000000000001011"), -- i=584
      ("01", "0000000000001001", "0000000000000010", "0000000000000111"), -- i=585
      ("10", "0000000000001001", "0000000000000010", "0000000000000000"), -- i=586
      ("11", "0000000000001001", "0000000000000010", "0000000000001011"), -- i=587
      ("00", "0000000000001001", "0000000000000011", "0000000000001100"), -- i=588
      ("01", "0000000000001001", "0000000000000011", "0000000000000110"), -- i=589
      ("10", "0000000000001001", "0000000000000011", "0000000000000001"), -- i=590
      ("11", "0000000000001001", "0000000000000011", "0000000000001011"), -- i=591
      ("00", "0000000000001001", "0000000000000100", "0000000000001101"), -- i=592
      ("01", "0000000000001001", "0000000000000100", "0000000000000101"), -- i=593
      ("10", "0000000000001001", "0000000000000100", "0000000000000000"), -- i=594
      ("11", "0000000000001001", "0000000000000100", "0000000000001101"), -- i=595
      ("00", "0000000000001001", "0000000000000101", "0000000000001110"), -- i=596
      ("01", "0000000000001001", "0000000000000101", "0000000000000100"), -- i=597
      ("10", "0000000000001001", "0000000000000101", "0000000000000001"), -- i=598
      ("11", "0000000000001001", "0000000000000101", "0000000000001101"), -- i=599
      ("00", "0000000000001001", "0000000000000110", "0000000000001111"), -- i=600
      ("01", "0000000000001001", "0000000000000110", "0000000000000011"), -- i=601
      ("10", "0000000000001001", "0000000000000110", "0000000000000000"), -- i=602
      ("11", "0000000000001001", "0000000000000110", "0000000000001111"), -- i=603
      ("00", "0000000000001001", "0000000000000111", "0000000000010000"), -- i=604
      ("01", "0000000000001001", "0000000000000111", "0000000000000010"), -- i=605
      ("10", "0000000000001001", "0000000000000111", "0000000000000001"), -- i=606
      ("11", "0000000000001001", "0000000000000111", "0000000000001111"), -- i=607
      ("00", "0000000000001001", "0000000000001000", "0000000000010001"), -- i=608
      ("01", "0000000000001001", "0000000000001000", "0000000000000001"), -- i=609
      ("10", "0000000000001001", "0000000000001000", "0000000000001000"), -- i=610
      ("11", "0000000000001001", "0000000000001000", "0000000000001001"), -- i=611
      ("00", "0000000000001001", "0000000000001001", "0000000000010010"), -- i=612
      ("01", "0000000000001001", "0000000000001001", "0000000000000000"), -- i=613
      ("10", "0000000000001001", "0000000000001001", "0000000000001001"), -- i=614
      ("11", "0000000000001001", "0000000000001001", "0000000000001001"), -- i=615
      ("00", "0000000000001001", "0000000000001010", "0000000000010011"), -- i=616
      ("01", "0000000000001001", "0000000000001010", "1111111111111111"), -- i=617
      ("10", "0000000000001001", "0000000000001010", "0000000000001000"), -- i=618
      ("11", "0000000000001001", "0000000000001010", "0000000000001011"), -- i=619
      ("00", "0000000000001001", "0000000000001011", "0000000000010100"), -- i=620
      ("01", "0000000000001001", "0000000000001011", "1111111111111110"), -- i=621
      ("10", "0000000000001001", "0000000000001011", "0000000000001001"), -- i=622
      ("11", "0000000000001001", "0000000000001011", "0000000000001011"), -- i=623
      ("00", "0000000000001001", "0000000000001100", "0000000000010101"), -- i=624
      ("01", "0000000000001001", "0000000000001100", "1111111111111101"), -- i=625
      ("10", "0000000000001001", "0000000000001100", "0000000000001000"), -- i=626
      ("11", "0000000000001001", "0000000000001100", "0000000000001101"), -- i=627
      ("00", "0000000000001001", "0000000000001101", "0000000000010110"), -- i=628
      ("01", "0000000000001001", "0000000000001101", "1111111111111100"), -- i=629
      ("10", "0000000000001001", "0000000000001101", "0000000000001001"), -- i=630
      ("11", "0000000000001001", "0000000000001101", "0000000000001101"), -- i=631
      ("00", "0000000000001001", "0000000000001110", "0000000000010111"), -- i=632
      ("01", "0000000000001001", "0000000000001110", "1111111111111011"), -- i=633
      ("10", "0000000000001001", "0000000000001110", "0000000000001000"), -- i=634
      ("11", "0000000000001001", "0000000000001110", "0000000000001111"), -- i=635
      ("00", "0000000000001001", "0000000000001111", "0000000000011000"), -- i=636
      ("01", "0000000000001001", "0000000000001111", "1111111111111010"), -- i=637
      ("10", "0000000000001001", "0000000000001111", "0000000000001001"), -- i=638
      ("11", "0000000000001001", "0000000000001111", "0000000000001111"), -- i=639
      ("00", "0000000000001010", "0000000000000000", "0000000000001010"), -- i=640
      ("01", "0000000000001010", "0000000000000000", "0000000000001010"), -- i=641
      ("10", "0000000000001010", "0000000000000000", "0000000000000000"), -- i=642
      ("11", "0000000000001010", "0000000000000000", "0000000000001010"), -- i=643
      ("00", "0000000000001010", "0000000000000001", "0000000000001011"), -- i=644
      ("01", "0000000000001010", "0000000000000001", "0000000000001001"), -- i=645
      ("10", "0000000000001010", "0000000000000001", "0000000000000000"), -- i=646
      ("11", "0000000000001010", "0000000000000001", "0000000000001011"), -- i=647
      ("00", "0000000000001010", "0000000000000010", "0000000000001100"), -- i=648
      ("01", "0000000000001010", "0000000000000010", "0000000000001000"), -- i=649
      ("10", "0000000000001010", "0000000000000010", "0000000000000010"), -- i=650
      ("11", "0000000000001010", "0000000000000010", "0000000000001010"), -- i=651
      ("00", "0000000000001010", "0000000000000011", "0000000000001101"), -- i=652
      ("01", "0000000000001010", "0000000000000011", "0000000000000111"), -- i=653
      ("10", "0000000000001010", "0000000000000011", "0000000000000010"), -- i=654
      ("11", "0000000000001010", "0000000000000011", "0000000000001011"), -- i=655
      ("00", "0000000000001010", "0000000000000100", "0000000000001110"), -- i=656
      ("01", "0000000000001010", "0000000000000100", "0000000000000110"), -- i=657
      ("10", "0000000000001010", "0000000000000100", "0000000000000000"), -- i=658
      ("11", "0000000000001010", "0000000000000100", "0000000000001110"), -- i=659
      ("00", "0000000000001010", "0000000000000101", "0000000000001111"), -- i=660
      ("01", "0000000000001010", "0000000000000101", "0000000000000101"), -- i=661
      ("10", "0000000000001010", "0000000000000101", "0000000000000000"), -- i=662
      ("11", "0000000000001010", "0000000000000101", "0000000000001111"), -- i=663
      ("00", "0000000000001010", "0000000000000110", "0000000000010000"), -- i=664
      ("01", "0000000000001010", "0000000000000110", "0000000000000100"), -- i=665
      ("10", "0000000000001010", "0000000000000110", "0000000000000010"), -- i=666
      ("11", "0000000000001010", "0000000000000110", "0000000000001110"), -- i=667
      ("00", "0000000000001010", "0000000000000111", "0000000000010001"), -- i=668
      ("01", "0000000000001010", "0000000000000111", "0000000000000011"), -- i=669
      ("10", "0000000000001010", "0000000000000111", "0000000000000010"), -- i=670
      ("11", "0000000000001010", "0000000000000111", "0000000000001111"), -- i=671
      ("00", "0000000000001010", "0000000000001000", "0000000000010010"), -- i=672
      ("01", "0000000000001010", "0000000000001000", "0000000000000010"), -- i=673
      ("10", "0000000000001010", "0000000000001000", "0000000000001000"), -- i=674
      ("11", "0000000000001010", "0000000000001000", "0000000000001010"), -- i=675
      ("00", "0000000000001010", "0000000000001001", "0000000000010011"), -- i=676
      ("01", "0000000000001010", "0000000000001001", "0000000000000001"), -- i=677
      ("10", "0000000000001010", "0000000000001001", "0000000000001000"), -- i=678
      ("11", "0000000000001010", "0000000000001001", "0000000000001011"), -- i=679
      ("00", "0000000000001010", "0000000000001010", "0000000000010100"), -- i=680
      ("01", "0000000000001010", "0000000000001010", "0000000000000000"), -- i=681
      ("10", "0000000000001010", "0000000000001010", "0000000000001010"), -- i=682
      ("11", "0000000000001010", "0000000000001010", "0000000000001010"), -- i=683
      ("00", "0000000000001010", "0000000000001011", "0000000000010101"), -- i=684
      ("01", "0000000000001010", "0000000000001011", "1111111111111111"), -- i=685
      ("10", "0000000000001010", "0000000000001011", "0000000000001010"), -- i=686
      ("11", "0000000000001010", "0000000000001011", "0000000000001011"), -- i=687
      ("00", "0000000000001010", "0000000000001100", "0000000000010110"), -- i=688
      ("01", "0000000000001010", "0000000000001100", "1111111111111110"), -- i=689
      ("10", "0000000000001010", "0000000000001100", "0000000000001000"), -- i=690
      ("11", "0000000000001010", "0000000000001100", "0000000000001110"), -- i=691
      ("00", "0000000000001010", "0000000000001101", "0000000000010111"), -- i=692
      ("01", "0000000000001010", "0000000000001101", "1111111111111101"), -- i=693
      ("10", "0000000000001010", "0000000000001101", "0000000000001000"), -- i=694
      ("11", "0000000000001010", "0000000000001101", "0000000000001111"), -- i=695
      ("00", "0000000000001010", "0000000000001110", "0000000000011000"), -- i=696
      ("01", "0000000000001010", "0000000000001110", "1111111111111100"), -- i=697
      ("10", "0000000000001010", "0000000000001110", "0000000000001010"), -- i=698
      ("11", "0000000000001010", "0000000000001110", "0000000000001110"), -- i=699
      ("00", "0000000000001010", "0000000000001111", "0000000000011001"), -- i=700
      ("01", "0000000000001010", "0000000000001111", "1111111111111011"), -- i=701
      ("10", "0000000000001010", "0000000000001111", "0000000000001010"), -- i=702
      ("11", "0000000000001010", "0000000000001111", "0000000000001111"), -- i=703
      ("00", "0000000000001011", "0000000000000000", "0000000000001011"), -- i=704
      ("01", "0000000000001011", "0000000000000000", "0000000000001011"), -- i=705
      ("10", "0000000000001011", "0000000000000000", "0000000000000000"), -- i=706
      ("11", "0000000000001011", "0000000000000000", "0000000000001011"), -- i=707
      ("00", "0000000000001011", "0000000000000001", "0000000000001100"), -- i=708
      ("01", "0000000000001011", "0000000000000001", "0000000000001010"), -- i=709
      ("10", "0000000000001011", "0000000000000001", "0000000000000001"), -- i=710
      ("11", "0000000000001011", "0000000000000001", "0000000000001011"), -- i=711
      ("00", "0000000000001011", "0000000000000010", "0000000000001101"), -- i=712
      ("01", "0000000000001011", "0000000000000010", "0000000000001001"), -- i=713
      ("10", "0000000000001011", "0000000000000010", "0000000000000010"), -- i=714
      ("11", "0000000000001011", "0000000000000010", "0000000000001011"), -- i=715
      ("00", "0000000000001011", "0000000000000011", "0000000000001110"), -- i=716
      ("01", "0000000000001011", "0000000000000011", "0000000000001000"), -- i=717
      ("10", "0000000000001011", "0000000000000011", "0000000000000011"), -- i=718
      ("11", "0000000000001011", "0000000000000011", "0000000000001011"), -- i=719
      ("00", "0000000000001011", "0000000000000100", "0000000000001111"), -- i=720
      ("01", "0000000000001011", "0000000000000100", "0000000000000111"), -- i=721
      ("10", "0000000000001011", "0000000000000100", "0000000000000000"), -- i=722
      ("11", "0000000000001011", "0000000000000100", "0000000000001111"), -- i=723
      ("00", "0000000000001011", "0000000000000101", "0000000000010000"), -- i=724
      ("01", "0000000000001011", "0000000000000101", "0000000000000110"), -- i=725
      ("10", "0000000000001011", "0000000000000101", "0000000000000001"), -- i=726
      ("11", "0000000000001011", "0000000000000101", "0000000000001111"), -- i=727
      ("00", "0000000000001011", "0000000000000110", "0000000000010001"), -- i=728
      ("01", "0000000000001011", "0000000000000110", "0000000000000101"), -- i=729
      ("10", "0000000000001011", "0000000000000110", "0000000000000010"), -- i=730
      ("11", "0000000000001011", "0000000000000110", "0000000000001111"), -- i=731
      ("00", "0000000000001011", "0000000000000111", "0000000000010010"), -- i=732
      ("01", "0000000000001011", "0000000000000111", "0000000000000100"), -- i=733
      ("10", "0000000000001011", "0000000000000111", "0000000000000011"), -- i=734
      ("11", "0000000000001011", "0000000000000111", "0000000000001111"), -- i=735
      ("00", "0000000000001011", "0000000000001000", "0000000000010011"), -- i=736
      ("01", "0000000000001011", "0000000000001000", "0000000000000011"), -- i=737
      ("10", "0000000000001011", "0000000000001000", "0000000000001000"), -- i=738
      ("11", "0000000000001011", "0000000000001000", "0000000000001011"), -- i=739
      ("00", "0000000000001011", "0000000000001001", "0000000000010100"), -- i=740
      ("01", "0000000000001011", "0000000000001001", "0000000000000010"), -- i=741
      ("10", "0000000000001011", "0000000000001001", "0000000000001001"), -- i=742
      ("11", "0000000000001011", "0000000000001001", "0000000000001011"), -- i=743
      ("00", "0000000000001011", "0000000000001010", "0000000000010101"), -- i=744
      ("01", "0000000000001011", "0000000000001010", "0000000000000001"), -- i=745
      ("10", "0000000000001011", "0000000000001010", "0000000000001010"), -- i=746
      ("11", "0000000000001011", "0000000000001010", "0000000000001011"), -- i=747
      ("00", "0000000000001011", "0000000000001011", "0000000000010110"), -- i=748
      ("01", "0000000000001011", "0000000000001011", "0000000000000000"), -- i=749
      ("10", "0000000000001011", "0000000000001011", "0000000000001011"), -- i=750
      ("11", "0000000000001011", "0000000000001011", "0000000000001011"), -- i=751
      ("00", "0000000000001011", "0000000000001100", "0000000000010111"), -- i=752
      ("01", "0000000000001011", "0000000000001100", "1111111111111111"), -- i=753
      ("10", "0000000000001011", "0000000000001100", "0000000000001000"), -- i=754
      ("11", "0000000000001011", "0000000000001100", "0000000000001111"), -- i=755
      ("00", "0000000000001011", "0000000000001101", "0000000000011000"), -- i=756
      ("01", "0000000000001011", "0000000000001101", "1111111111111110"), -- i=757
      ("10", "0000000000001011", "0000000000001101", "0000000000001001"), -- i=758
      ("11", "0000000000001011", "0000000000001101", "0000000000001111"), -- i=759
      ("00", "0000000000001011", "0000000000001110", "0000000000011001"), -- i=760
      ("01", "0000000000001011", "0000000000001110", "1111111111111101"), -- i=761
      ("10", "0000000000001011", "0000000000001110", "0000000000001010"), -- i=762
      ("11", "0000000000001011", "0000000000001110", "0000000000001111"), -- i=763
      ("00", "0000000000001011", "0000000000001111", "0000000000011010"), -- i=764
      ("01", "0000000000001011", "0000000000001111", "1111111111111100"), -- i=765
      ("10", "0000000000001011", "0000000000001111", "0000000000001011"), -- i=766
      ("11", "0000000000001011", "0000000000001111", "0000000000001111"), -- i=767
      ("00", "0000000000001100", "0000000000000000", "0000000000001100"), -- i=768
      ("01", "0000000000001100", "0000000000000000", "0000000000001100"), -- i=769
      ("10", "0000000000001100", "0000000000000000", "0000000000000000"), -- i=770
      ("11", "0000000000001100", "0000000000000000", "0000000000001100"), -- i=771
      ("00", "0000000000001100", "0000000000000001", "0000000000001101"), -- i=772
      ("01", "0000000000001100", "0000000000000001", "0000000000001011"), -- i=773
      ("10", "0000000000001100", "0000000000000001", "0000000000000000"), -- i=774
      ("11", "0000000000001100", "0000000000000001", "0000000000001101"), -- i=775
      ("00", "0000000000001100", "0000000000000010", "0000000000001110"), -- i=776
      ("01", "0000000000001100", "0000000000000010", "0000000000001010"), -- i=777
      ("10", "0000000000001100", "0000000000000010", "0000000000000000"), -- i=778
      ("11", "0000000000001100", "0000000000000010", "0000000000001110"), -- i=779
      ("00", "0000000000001100", "0000000000000011", "0000000000001111"), -- i=780
      ("01", "0000000000001100", "0000000000000011", "0000000000001001"), -- i=781
      ("10", "0000000000001100", "0000000000000011", "0000000000000000"), -- i=782
      ("11", "0000000000001100", "0000000000000011", "0000000000001111"), -- i=783
      ("00", "0000000000001100", "0000000000000100", "0000000000010000"), -- i=784
      ("01", "0000000000001100", "0000000000000100", "0000000000001000"), -- i=785
      ("10", "0000000000001100", "0000000000000100", "0000000000000100"), -- i=786
      ("11", "0000000000001100", "0000000000000100", "0000000000001100"), -- i=787
      ("00", "0000000000001100", "0000000000000101", "0000000000010001"), -- i=788
      ("01", "0000000000001100", "0000000000000101", "0000000000000111"), -- i=789
      ("10", "0000000000001100", "0000000000000101", "0000000000000100"), -- i=790
      ("11", "0000000000001100", "0000000000000101", "0000000000001101"), -- i=791
      ("00", "0000000000001100", "0000000000000110", "0000000000010010"), -- i=792
      ("01", "0000000000001100", "0000000000000110", "0000000000000110"), -- i=793
      ("10", "0000000000001100", "0000000000000110", "0000000000000100"), -- i=794
      ("11", "0000000000001100", "0000000000000110", "0000000000001110"), -- i=795
      ("00", "0000000000001100", "0000000000000111", "0000000000010011"), -- i=796
      ("01", "0000000000001100", "0000000000000111", "0000000000000101"), -- i=797
      ("10", "0000000000001100", "0000000000000111", "0000000000000100"), -- i=798
      ("11", "0000000000001100", "0000000000000111", "0000000000001111"), -- i=799
      ("00", "0000000000001100", "0000000000001000", "0000000000010100"), -- i=800
      ("01", "0000000000001100", "0000000000001000", "0000000000000100"), -- i=801
      ("10", "0000000000001100", "0000000000001000", "0000000000001000"), -- i=802
      ("11", "0000000000001100", "0000000000001000", "0000000000001100"), -- i=803
      ("00", "0000000000001100", "0000000000001001", "0000000000010101"), -- i=804
      ("01", "0000000000001100", "0000000000001001", "0000000000000011"), -- i=805
      ("10", "0000000000001100", "0000000000001001", "0000000000001000"), -- i=806
      ("11", "0000000000001100", "0000000000001001", "0000000000001101"), -- i=807
      ("00", "0000000000001100", "0000000000001010", "0000000000010110"), -- i=808
      ("01", "0000000000001100", "0000000000001010", "0000000000000010"), -- i=809
      ("10", "0000000000001100", "0000000000001010", "0000000000001000"), -- i=810
      ("11", "0000000000001100", "0000000000001010", "0000000000001110"), -- i=811
      ("00", "0000000000001100", "0000000000001011", "0000000000010111"), -- i=812
      ("01", "0000000000001100", "0000000000001011", "0000000000000001"), -- i=813
      ("10", "0000000000001100", "0000000000001011", "0000000000001000"), -- i=814
      ("11", "0000000000001100", "0000000000001011", "0000000000001111"), -- i=815
      ("00", "0000000000001100", "0000000000001100", "0000000000011000"), -- i=816
      ("01", "0000000000001100", "0000000000001100", "0000000000000000"), -- i=817
      ("10", "0000000000001100", "0000000000001100", "0000000000001100"), -- i=818
      ("11", "0000000000001100", "0000000000001100", "0000000000001100"), -- i=819
      ("00", "0000000000001100", "0000000000001101", "0000000000011001"), -- i=820
      ("01", "0000000000001100", "0000000000001101", "1111111111111111"), -- i=821
      ("10", "0000000000001100", "0000000000001101", "0000000000001100"), -- i=822
      ("11", "0000000000001100", "0000000000001101", "0000000000001101"), -- i=823
      ("00", "0000000000001100", "0000000000001110", "0000000000011010"), -- i=824
      ("01", "0000000000001100", "0000000000001110", "1111111111111110"), -- i=825
      ("10", "0000000000001100", "0000000000001110", "0000000000001100"), -- i=826
      ("11", "0000000000001100", "0000000000001110", "0000000000001110"), -- i=827
      ("00", "0000000000001100", "0000000000001111", "0000000000011011"), -- i=828
      ("01", "0000000000001100", "0000000000001111", "1111111111111101"), -- i=829
      ("10", "0000000000001100", "0000000000001111", "0000000000001100"), -- i=830
      ("11", "0000000000001100", "0000000000001111", "0000000000001111"), -- i=831
      ("00", "0000000000001101", "0000000000000000", "0000000000001101"), -- i=832
      ("01", "0000000000001101", "0000000000000000", "0000000000001101"), -- i=833
      ("10", "0000000000001101", "0000000000000000", "0000000000000000"), -- i=834
      ("11", "0000000000001101", "0000000000000000", "0000000000001101"), -- i=835
      ("00", "0000000000001101", "0000000000000001", "0000000000001110"), -- i=836
      ("01", "0000000000001101", "0000000000000001", "0000000000001100"), -- i=837
      ("10", "0000000000001101", "0000000000000001", "0000000000000001"), -- i=838
      ("11", "0000000000001101", "0000000000000001", "0000000000001101"), -- i=839
      ("00", "0000000000001101", "0000000000000010", "0000000000001111"), -- i=840
      ("01", "0000000000001101", "0000000000000010", "0000000000001011"), -- i=841
      ("10", "0000000000001101", "0000000000000010", "0000000000000000"), -- i=842
      ("11", "0000000000001101", "0000000000000010", "0000000000001111"), -- i=843
      ("00", "0000000000001101", "0000000000000011", "0000000000010000"), -- i=844
      ("01", "0000000000001101", "0000000000000011", "0000000000001010"), -- i=845
      ("10", "0000000000001101", "0000000000000011", "0000000000000001"), -- i=846
      ("11", "0000000000001101", "0000000000000011", "0000000000001111"), -- i=847
      ("00", "0000000000001101", "0000000000000100", "0000000000010001"), -- i=848
      ("01", "0000000000001101", "0000000000000100", "0000000000001001"), -- i=849
      ("10", "0000000000001101", "0000000000000100", "0000000000000100"), -- i=850
      ("11", "0000000000001101", "0000000000000100", "0000000000001101"), -- i=851
      ("00", "0000000000001101", "0000000000000101", "0000000000010010"), -- i=852
      ("01", "0000000000001101", "0000000000000101", "0000000000001000"), -- i=853
      ("10", "0000000000001101", "0000000000000101", "0000000000000101"), -- i=854
      ("11", "0000000000001101", "0000000000000101", "0000000000001101"), -- i=855
      ("00", "0000000000001101", "0000000000000110", "0000000000010011"), -- i=856
      ("01", "0000000000001101", "0000000000000110", "0000000000000111"), -- i=857
      ("10", "0000000000001101", "0000000000000110", "0000000000000100"), -- i=858
      ("11", "0000000000001101", "0000000000000110", "0000000000001111"), -- i=859
      ("00", "0000000000001101", "0000000000000111", "0000000000010100"), -- i=860
      ("01", "0000000000001101", "0000000000000111", "0000000000000110"), -- i=861
      ("10", "0000000000001101", "0000000000000111", "0000000000000101"), -- i=862
      ("11", "0000000000001101", "0000000000000111", "0000000000001111"), -- i=863
      ("00", "0000000000001101", "0000000000001000", "0000000000010101"), -- i=864
      ("01", "0000000000001101", "0000000000001000", "0000000000000101"), -- i=865
      ("10", "0000000000001101", "0000000000001000", "0000000000001000"), -- i=866
      ("11", "0000000000001101", "0000000000001000", "0000000000001101"), -- i=867
      ("00", "0000000000001101", "0000000000001001", "0000000000010110"), -- i=868
      ("01", "0000000000001101", "0000000000001001", "0000000000000100"), -- i=869
      ("10", "0000000000001101", "0000000000001001", "0000000000001001"), -- i=870
      ("11", "0000000000001101", "0000000000001001", "0000000000001101"), -- i=871
      ("00", "0000000000001101", "0000000000001010", "0000000000010111"), -- i=872
      ("01", "0000000000001101", "0000000000001010", "0000000000000011"), -- i=873
      ("10", "0000000000001101", "0000000000001010", "0000000000001000"), -- i=874
      ("11", "0000000000001101", "0000000000001010", "0000000000001111"), -- i=875
      ("00", "0000000000001101", "0000000000001011", "0000000000011000"), -- i=876
      ("01", "0000000000001101", "0000000000001011", "0000000000000010"), -- i=877
      ("10", "0000000000001101", "0000000000001011", "0000000000001001"), -- i=878
      ("11", "0000000000001101", "0000000000001011", "0000000000001111"), -- i=879
      ("00", "0000000000001101", "0000000000001100", "0000000000011001"), -- i=880
      ("01", "0000000000001101", "0000000000001100", "0000000000000001"), -- i=881
      ("10", "0000000000001101", "0000000000001100", "0000000000001100"), -- i=882
      ("11", "0000000000001101", "0000000000001100", "0000000000001101"), -- i=883
      ("00", "0000000000001101", "0000000000001101", "0000000000011010"), -- i=884
      ("01", "0000000000001101", "0000000000001101", "0000000000000000"), -- i=885
      ("10", "0000000000001101", "0000000000001101", "0000000000001101"), -- i=886
      ("11", "0000000000001101", "0000000000001101", "0000000000001101"), -- i=887
      ("00", "0000000000001101", "0000000000001110", "0000000000011011"), -- i=888
      ("01", "0000000000001101", "0000000000001110", "1111111111111111"), -- i=889
      ("10", "0000000000001101", "0000000000001110", "0000000000001100"), -- i=890
      ("11", "0000000000001101", "0000000000001110", "0000000000001111"), -- i=891
      ("00", "0000000000001101", "0000000000001111", "0000000000011100"), -- i=892
      ("01", "0000000000001101", "0000000000001111", "1111111111111110"), -- i=893
      ("10", "0000000000001101", "0000000000001111", "0000000000001101"), -- i=894
      ("11", "0000000000001101", "0000000000001111", "0000000000001111"), -- i=895
      ("00", "0000000000001110", "0000000000000000", "0000000000001110"), -- i=896
      ("01", "0000000000001110", "0000000000000000", "0000000000001110"), -- i=897
      ("10", "0000000000001110", "0000000000000000", "0000000000000000"), -- i=898
      ("11", "0000000000001110", "0000000000000000", "0000000000001110"), -- i=899
      ("00", "0000000000001110", "0000000000000001", "0000000000001111"), -- i=900
      ("01", "0000000000001110", "0000000000000001", "0000000000001101"), -- i=901
      ("10", "0000000000001110", "0000000000000001", "0000000000000000"), -- i=902
      ("11", "0000000000001110", "0000000000000001", "0000000000001111"), -- i=903
      ("00", "0000000000001110", "0000000000000010", "0000000000010000"), -- i=904
      ("01", "0000000000001110", "0000000000000010", "0000000000001100"), -- i=905
      ("10", "0000000000001110", "0000000000000010", "0000000000000010"), -- i=906
      ("11", "0000000000001110", "0000000000000010", "0000000000001110"), -- i=907
      ("00", "0000000000001110", "0000000000000011", "0000000000010001"), -- i=908
      ("01", "0000000000001110", "0000000000000011", "0000000000001011"), -- i=909
      ("10", "0000000000001110", "0000000000000011", "0000000000000010"), -- i=910
      ("11", "0000000000001110", "0000000000000011", "0000000000001111"), -- i=911
      ("00", "0000000000001110", "0000000000000100", "0000000000010010"), -- i=912
      ("01", "0000000000001110", "0000000000000100", "0000000000001010"), -- i=913
      ("10", "0000000000001110", "0000000000000100", "0000000000000100"), -- i=914
      ("11", "0000000000001110", "0000000000000100", "0000000000001110"), -- i=915
      ("00", "0000000000001110", "0000000000000101", "0000000000010011"), -- i=916
      ("01", "0000000000001110", "0000000000000101", "0000000000001001"), -- i=917
      ("10", "0000000000001110", "0000000000000101", "0000000000000100"), -- i=918
      ("11", "0000000000001110", "0000000000000101", "0000000000001111"), -- i=919
      ("00", "0000000000001110", "0000000000000110", "0000000000010100"), -- i=920
      ("01", "0000000000001110", "0000000000000110", "0000000000001000"), -- i=921
      ("10", "0000000000001110", "0000000000000110", "0000000000000110"), -- i=922
      ("11", "0000000000001110", "0000000000000110", "0000000000001110"), -- i=923
      ("00", "0000000000001110", "0000000000000111", "0000000000010101"), -- i=924
      ("01", "0000000000001110", "0000000000000111", "0000000000000111"), -- i=925
      ("10", "0000000000001110", "0000000000000111", "0000000000000110"), -- i=926
      ("11", "0000000000001110", "0000000000000111", "0000000000001111"), -- i=927
      ("00", "0000000000001110", "0000000000001000", "0000000000010110"), -- i=928
      ("01", "0000000000001110", "0000000000001000", "0000000000000110"), -- i=929
      ("10", "0000000000001110", "0000000000001000", "0000000000001000"), -- i=930
      ("11", "0000000000001110", "0000000000001000", "0000000000001110"), -- i=931
      ("00", "0000000000001110", "0000000000001001", "0000000000010111"), -- i=932
      ("01", "0000000000001110", "0000000000001001", "0000000000000101"), -- i=933
      ("10", "0000000000001110", "0000000000001001", "0000000000001000"), -- i=934
      ("11", "0000000000001110", "0000000000001001", "0000000000001111"), -- i=935
      ("00", "0000000000001110", "0000000000001010", "0000000000011000"), -- i=936
      ("01", "0000000000001110", "0000000000001010", "0000000000000100"), -- i=937
      ("10", "0000000000001110", "0000000000001010", "0000000000001010"), -- i=938
      ("11", "0000000000001110", "0000000000001010", "0000000000001110"), -- i=939
      ("00", "0000000000001110", "0000000000001011", "0000000000011001"), -- i=940
      ("01", "0000000000001110", "0000000000001011", "0000000000000011"), -- i=941
      ("10", "0000000000001110", "0000000000001011", "0000000000001010"), -- i=942
      ("11", "0000000000001110", "0000000000001011", "0000000000001111"), -- i=943
      ("00", "0000000000001110", "0000000000001100", "0000000000011010"), -- i=944
      ("01", "0000000000001110", "0000000000001100", "0000000000000010"), -- i=945
      ("10", "0000000000001110", "0000000000001100", "0000000000001100"), -- i=946
      ("11", "0000000000001110", "0000000000001100", "0000000000001110"), -- i=947
      ("00", "0000000000001110", "0000000000001101", "0000000000011011"), -- i=948
      ("01", "0000000000001110", "0000000000001101", "0000000000000001"), -- i=949
      ("10", "0000000000001110", "0000000000001101", "0000000000001100"), -- i=950
      ("11", "0000000000001110", "0000000000001101", "0000000000001111"), -- i=951
      ("00", "0000000000001110", "0000000000001110", "0000000000011100"), -- i=952
      ("01", "0000000000001110", "0000000000001110", "0000000000000000"), -- i=953
      ("10", "0000000000001110", "0000000000001110", "0000000000001110"), -- i=954
      ("11", "0000000000001110", "0000000000001110", "0000000000001110"), -- i=955
      ("00", "0000000000001110", "0000000000001111", "0000000000011101"), -- i=956
      ("01", "0000000000001110", "0000000000001111", "1111111111111111"), -- i=957
      ("10", "0000000000001110", "0000000000001111", "0000000000001110"), -- i=958
      ("11", "0000000000001110", "0000000000001111", "0000000000001111"), -- i=959
      ("00", "0000000000001111", "0000000000000000", "0000000000001111"), -- i=960
      ("01", "0000000000001111", "0000000000000000", "0000000000001111"), -- i=961
      ("10", "0000000000001111", "0000000000000000", "0000000000000000"), -- i=962
      ("11", "0000000000001111", "0000000000000000", "0000000000001111"), -- i=963
      ("00", "0000000000001111", "0000000000000001", "0000000000010000"), -- i=964
      ("01", "0000000000001111", "0000000000000001", "0000000000001110"), -- i=965
      ("10", "0000000000001111", "0000000000000001", "0000000000000001"), -- i=966
      ("11", "0000000000001111", "0000000000000001", "0000000000001111"), -- i=967
      ("00", "0000000000001111", "0000000000000010", "0000000000010001"), -- i=968
      ("01", "0000000000001111", "0000000000000010", "0000000000001101"), -- i=969
      ("10", "0000000000001111", "0000000000000010", "0000000000000010"), -- i=970
      ("11", "0000000000001111", "0000000000000010", "0000000000001111"), -- i=971
      ("00", "0000000000001111", "0000000000000011", "0000000000010010"), -- i=972
      ("01", "0000000000001111", "0000000000000011", "0000000000001100"), -- i=973
      ("10", "0000000000001111", "0000000000000011", "0000000000000011"), -- i=974
      ("11", "0000000000001111", "0000000000000011", "0000000000001111"), -- i=975
      ("00", "0000000000001111", "0000000000000100", "0000000000010011"), -- i=976
      ("01", "0000000000001111", "0000000000000100", "0000000000001011"), -- i=977
      ("10", "0000000000001111", "0000000000000100", "0000000000000100"), -- i=978
      ("11", "0000000000001111", "0000000000000100", "0000000000001111"), -- i=979
      ("00", "0000000000001111", "0000000000000101", "0000000000010100"), -- i=980
      ("01", "0000000000001111", "0000000000000101", "0000000000001010"), -- i=981
      ("10", "0000000000001111", "0000000000000101", "0000000000000101"), -- i=982
      ("11", "0000000000001111", "0000000000000101", "0000000000001111"), -- i=983
      ("00", "0000000000001111", "0000000000000110", "0000000000010101"), -- i=984
      ("01", "0000000000001111", "0000000000000110", "0000000000001001"), -- i=985
      ("10", "0000000000001111", "0000000000000110", "0000000000000110"), -- i=986
      ("11", "0000000000001111", "0000000000000110", "0000000000001111"), -- i=987
      ("00", "0000000000001111", "0000000000000111", "0000000000010110"), -- i=988
      ("01", "0000000000001111", "0000000000000111", "0000000000001000"), -- i=989
      ("10", "0000000000001111", "0000000000000111", "0000000000000111"), -- i=990
      ("11", "0000000000001111", "0000000000000111", "0000000000001111"), -- i=991
      ("00", "0000000000001111", "0000000000001000", "0000000000010111"), -- i=992
      ("01", "0000000000001111", "0000000000001000", "0000000000000111"), -- i=993
      ("10", "0000000000001111", "0000000000001000", "0000000000001000"), -- i=994
      ("11", "0000000000001111", "0000000000001000", "0000000000001111"), -- i=995
      ("00", "0000000000001111", "0000000000001001", "0000000000011000"), -- i=996
      ("01", "0000000000001111", "0000000000001001", "0000000000000110"), -- i=997
      ("10", "0000000000001111", "0000000000001001", "0000000000001001"), -- i=998
      ("11", "0000000000001111", "0000000000001001", "0000000000001111"), -- i=999
      ("00", "0000000000001111", "0000000000001010", "0000000000011001"), -- i=1000
      ("01", "0000000000001111", "0000000000001010", "0000000000000101"), -- i=1001
      ("10", "0000000000001111", "0000000000001010", "0000000000001010"), -- i=1002
      ("11", "0000000000001111", "0000000000001010", "0000000000001111"), -- i=1003
      ("00", "0000000000001111", "0000000000001011", "0000000000011010"), -- i=1004
      ("01", "0000000000001111", "0000000000001011", "0000000000000100"), -- i=1005
      ("10", "0000000000001111", "0000000000001011", "0000000000001011"), -- i=1006
      ("11", "0000000000001111", "0000000000001011", "0000000000001111"), -- i=1007
      ("00", "0000000000001111", "0000000000001100", "0000000000011011"), -- i=1008
      ("01", "0000000000001111", "0000000000001100", "0000000000000011"), -- i=1009
      ("10", "0000000000001111", "0000000000001100", "0000000000001100"), -- i=1010
      ("11", "0000000000001111", "0000000000001100", "0000000000001111"), -- i=1011
      ("00", "0000000000001111", "0000000000001101", "0000000000011100"), -- i=1012
      ("01", "0000000000001111", "0000000000001101", "0000000000000010"), -- i=1013
      ("10", "0000000000001111", "0000000000001101", "0000000000001101"), -- i=1014
      ("11", "0000000000001111", "0000000000001101", "0000000000001111"), -- i=1015
      ("00", "0000000000001111", "0000000000001110", "0000000000011101"), -- i=1016
      ("01", "0000000000001111", "0000000000001110", "0000000000000001"), -- i=1017
      ("10", "0000000000001111", "0000000000001110", "0000000000001110"), -- i=1018
      ("11", "0000000000001111", "0000000000001110", "0000000000001111"), -- i=1019
      ("00", "0000000000001111", "0000000000001111", "0000000000011110"), -- i=1020
      ("01", "0000000000001111", "0000000000001111", "0000000000000000"), -- i=1021
      ("10", "0000000000001111", "0000000000001111", "0000000000001111"), -- i=1022
      ("11", "0000000000001111", "0000000000001111", "0000000000001111"), -- i=1023
      ("00", "1101111011101000", "0111000010100000", "0100111110001000"), -- i=1024
      ("01", "1101111011101000", "0111000010100000", "0110111001001000"), -- i=1025
      ("10", "1101111011101000", "0111000010100000", "0101000010100000"), -- i=1026
      ("11", "1101111011101000", "0111000010100000", "1111111011101000"), -- i=1027
      ("00", "1001011111010011", "0010010001101000", "1011110000111011"), -- i=1028
      ("01", "1001011111010011", "0010010001101000", "0111001101101011"), -- i=1029
      ("10", "1001011111010011", "0010010001101000", "0000010001000000"), -- i=1030
      ("11", "1001011111010011", "0010010001101000", "1011011111111011"), -- i=1031
      ("00", "1000000101100101", "0111111010110010", "0000000000010111"), -- i=1032
      ("01", "1000000101100101", "0111111010110010", "0000001010110011"), -- i=1033
      ("10", "1000000101100101", "0111111010110010", "0000000000100000"), -- i=1034
      ("11", "1000000101100101", "0111111010110010", "1111111111110111"), -- i=1035
      ("00", "1001100100110011", "0011100000111010", "1101000101101101"), -- i=1036
      ("01", "1001100100110011", "0011100000111010", "0110000011111001"), -- i=1037
      ("10", "1001100100110011", "0011100000111010", "0001100000110010"), -- i=1038
      ("11", "1001100100110011", "0011100000111010", "1011100100111011"), -- i=1039
      ("00", "1101001000100101", "0011100001001111", "0000101001110100"), -- i=1040
      ("01", "1101001000100101", "0011100001001111", "1001100111010110"), -- i=1041
      ("10", "1101001000100101", "0011100001001111", "0001000000000101"), -- i=1042
      ("11", "1101001000100101", "0011100001001111", "1111101001101111"), -- i=1043
      ("00", "0001000011110100", "1111000100000000", "0000000111110100"), -- i=1044
      ("01", "0001000011110100", "1111000100000000", "0001111111110100"), -- i=1045
      ("10", "0001000011110100", "1111000100000000", "0001000000000000"), -- i=1046
      ("11", "0001000011110100", "1111000100000000", "1111000111110100"), -- i=1047
      ("00", "0110110001111010", "0011011001111100", "1010001011110110"), -- i=1048
      ("01", "0110110001111010", "0011011001111100", "0011010111111110"), -- i=1049
      ("10", "0110110001111010", "0011011001111100", "0010010001111000"), -- i=1050
      ("11", "0110110001111010", "0011011001111100", "0111111001111110"), -- i=1051
      ("00", "1110000110000100", "1001101011001000", "0111110001001100"), -- i=1052
      ("01", "1110000110000100", "1001101011001000", "0100011010111100"), -- i=1053
      ("10", "1110000110000100", "1001101011001000", "1000000010000000"), -- i=1054
      ("11", "1110000110000100", "1001101011001000", "1111101111001100"), -- i=1055
      ("00", "0111001100101011", "1111100001001000", "0110101101110011"), -- i=1056
      ("01", "0111001100101011", "1111100001001000", "0111101011100011"), -- i=1057
      ("10", "0111001100101011", "1111100001001000", "0111000000001000"), -- i=1058
      ("11", "0111001100101011", "1111100001001000", "1111101101101011"), -- i=1059
      ("00", "1110011000110011", "1100011111110110", "1010111000101001"), -- i=1060
      ("01", "1110011000110011", "1100011111110110", "0001111000111101"), -- i=1061
      ("10", "1110011000110011", "1100011111110110", "1100011000110010"), -- i=1062
      ("11", "1110011000110011", "1100011111110110", "1110011111110111"), -- i=1063
      ("00", "1001110110101001", "1111101000011110", "1001011111000111"), -- i=1064
      ("01", "1001110110101001", "1111101000011110", "1010001110001011"), -- i=1065
      ("10", "1001110110101001", "1111101000011110", "1001100000001000"), -- i=1066
      ("11", "1001110110101001", "1111101000011110", "1111111110111111"), -- i=1067
      ("00", "0110000101011010", "0101010111111011", "1011011101010101"), -- i=1068
      ("01", "0110000101011010", "0101010111111011", "0000101101011111"), -- i=1069
      ("10", "0110000101011010", "0101010111111011", "0100000101011010"), -- i=1070
      ("11", "0110000101011010", "0101010111111011", "0111010111111011"), -- i=1071
      ("00", "0010000111101010", "0110010001000101", "1000011000101111"), -- i=1072
      ("01", "0010000111101010", "0110010001000101", "1011110110100101"), -- i=1073
      ("10", "0010000111101010", "0110010001000101", "0010000001000000"), -- i=1074
      ("11", "0010000111101010", "0110010001000101", "0110010111101111"), -- i=1075
      ("00", "1101001010010000", "1100111001000001", "1010000011010001"), -- i=1076
      ("01", "1101001010010000", "1100111001000001", "0000010001001111"), -- i=1077
      ("10", "1101001010010000", "1100111001000001", "1100001000000000"), -- i=1078
      ("11", "1101001010010000", "1100111001000001", "1101111011010001"), -- i=1079
      ("00", "1011010000010000", "0000110101110111", "1100000110000111"), -- i=1080
      ("01", "1011010000010000", "0000110101110111", "1010011010011001"), -- i=1081
      ("10", "1011010000010000", "0000110101110111", "0000010000010000"), -- i=1082
      ("11", "1011010000010000", "0000110101110111", "1011110101110111"), -- i=1083
      ("00", "1000011111001000", "1010001010111101", "0010101010000101"), -- i=1084
      ("01", "1000011111001000", "1010001010111101", "1110010100001011"), -- i=1085
      ("10", "1000011111001000", "1010001010111101", "1000001010001000"), -- i=1086
      ("11", "1000011111001000", "1010001010111101", "1010011111111101"), -- i=1087
      ("00", "0000001001101011", "1001110101111011", "1001111111100110"), -- i=1088
      ("01", "0000001001101011", "1001110101111011", "0110010011110000"), -- i=1089
      ("10", "0000001001101011", "1001110101111011", "0000000001101011"), -- i=1090
      ("11", "0000001001101011", "1001110101111011", "1001111101111011"), -- i=1091
      ("00", "1111110101111010", "1000100011010001", "1000011001001011"), -- i=1092
      ("01", "1111110101111010", "1000100011010001", "0111010010101001"), -- i=1093
      ("10", "1111110101111010", "1000100011010001", "1000100001010000"), -- i=1094
      ("11", "1111110101111010", "1000100011010001", "1111110111111011"), -- i=1095
      ("00", "1010100101110111", "0101001100100000", "1111110010010111"), -- i=1096
      ("01", "1010100101110111", "0101001100100000", "0101011001010111"), -- i=1097
      ("10", "1010100101110111", "0101001100100000", "0000000100100000"), -- i=1098
      ("11", "1010100101110111", "0101001100100000", "1111101101110111"), -- i=1099
      ("00", "1100101100101010", "0010000001100000", "1110101110001010"), -- i=1100
      ("01", "1100101100101010", "0010000001100000", "1010101011001010"), -- i=1101
      ("10", "1100101100101010", "0010000001100000", "0000000000100000"), -- i=1102
      ("11", "1100101100101010", "0010000001100000", "1110101101101010"), -- i=1103
      ("00", "1001100011101101", "0101000000100001", "1110100100001110"), -- i=1104
      ("01", "1001100011101101", "0101000000100001", "0100100011001100"), -- i=1105
      ("10", "1001100011101101", "0101000000100001", "0001000000100001"), -- i=1106
      ("11", "1001100011101101", "0101000000100001", "1101100011101101"), -- i=1107
      ("00", "0110101011100000", "0010100001001100", "1001001100101100"), -- i=1108
      ("01", "0110101011100000", "0010100001001100", "0100001010010100"), -- i=1109
      ("10", "0110101011100000", "0010100001001100", "0010100001000000"), -- i=1110
      ("11", "0110101011100000", "0010100001001100", "0110101011101100"), -- i=1111
      ("00", "0100100000001100", "0101010010101101", "1001110010111001"), -- i=1112
      ("01", "0100100000001100", "0101010010101101", "1111001101011111"), -- i=1113
      ("10", "0100100000001100", "0101010010101101", "0100000000001100"), -- i=1114
      ("11", "0100100000001100", "0101010010101101", "0101110010101101"), -- i=1115
      ("00", "1010001101111110", "1011110010111000", "0110000000110110"), -- i=1116
      ("01", "1010001101111110", "1011110010111000", "1110011011000110"), -- i=1117
      ("10", "1010001101111110", "1011110010111000", "1010000000111000"), -- i=1118
      ("11", "1010001101111110", "1011110010111000", "1011111111111110"), -- i=1119
      ("00", "1110010010010111", "1000001110110000", "0110100001000111"), -- i=1120
      ("01", "1110010010010111", "1000001110110000", "0110000011100111"), -- i=1121
      ("10", "1110010010010111", "1000001110110000", "1000000010010000"), -- i=1122
      ("11", "1110010010010111", "1000001110110000", "1110011110110111"), -- i=1123
      ("00", "1011111100000001", "0111111011000011", "0011110111000100"), -- i=1124
      ("01", "1011111100000001", "0111111011000011", "0100000000111110"), -- i=1125
      ("10", "1011111100000001", "0111111011000011", "0011111000000001"), -- i=1126
      ("11", "1011111100000001", "0111111011000011", "1111111111000011"), -- i=1127
      ("00", "1101110101001000", "0010000000100000", "1111110101101000"), -- i=1128
      ("01", "1101110101001000", "0010000000100000", "1011110100101000"), -- i=1129
      ("10", "1101110101001000", "0010000000100000", "0000000000000000"), -- i=1130
      ("11", "1101110101001000", "0010000000100000", "1111110101101000"), -- i=1131
      ("00", "1111111100000100", "0001000010100101", "0000111110101001"), -- i=1132
      ("01", "1111111100000100", "0001000010100101", "1110111001011111"), -- i=1133
      ("10", "1111111100000100", "0001000010100101", "0001000000000100"), -- i=1134
      ("11", "1111111100000100", "0001000010100101", "1111111110100101"), -- i=1135
      ("00", "1100010110110110", "0011001011001110", "1111100010000100"), -- i=1136
      ("01", "1100010110110110", "0011001011001110", "1001001011101000"), -- i=1137
      ("10", "1100010110110110", "0011001011001110", "0000000010000110"), -- i=1138
      ("11", "1100010110110110", "0011001011001110", "1111011111111110"), -- i=1139
      ("00", "1111001100101001", "0000010001010011", "1111011101111100"), -- i=1140
      ("01", "1111001100101001", "0000010001010011", "1110111011010110"), -- i=1141
      ("10", "1111001100101001", "0000010001010011", "0000000000000001"), -- i=1142
      ("11", "1111001100101001", "0000010001010011", "1111011101111011"), -- i=1143
      ("00", "1001011011010011", "1010111110011010", "0100011001101101"), -- i=1144
      ("01", "1001011011010011", "1010111110011010", "1110011100111001"), -- i=1145
      ("10", "1001011011010011", "1010111110011010", "1000011010010010"), -- i=1146
      ("11", "1001011011010011", "1010111110011010", "1011111111011011"), -- i=1147
      ("00", "0110111000111101", "0011011000010110", "1010010001010011"), -- i=1148
      ("01", "0110111000111101", "0011011000010110", "0011100000100111"), -- i=1149
      ("10", "0110111000111101", "0011011000010110", "0010011000010100"), -- i=1150
      ("11", "0110111000111101", "0011011000010110", "0111111000111111"), -- i=1151
      ("00", "1011110010011011", "1111111111111001", "1011110010010100"), -- i=1152
      ("01", "1011110010011011", "1111111111111001", "1011110010100010"), -- i=1153
      ("10", "1011110010011011", "1111111111111001", "1011110010011001"), -- i=1154
      ("11", "1011110010011011", "1111111111111001", "1111111111111011"), -- i=1155
      ("00", "1101100000101111", "1000111111000010", "0110011111110001"), -- i=1156
      ("01", "1101100000101111", "1000111111000010", "0100100001101101"), -- i=1157
      ("10", "1101100000101111", "1000111111000010", "1000100000000010"), -- i=1158
      ("11", "1101100000101111", "1000111111000010", "1101111111101111"), -- i=1159
      ("00", "0011011010001100", "1101000000110100", "0000011011000000"), -- i=1160
      ("01", "0011011010001100", "1101000000110100", "0110011001011000"), -- i=1161
      ("10", "0011011010001100", "1101000000110100", "0001000000000100"), -- i=1162
      ("11", "0011011010001100", "1101000000110100", "1111011010111100"), -- i=1163
      ("00", "1000010000111000", "0101110001110110", "1110000010101110"), -- i=1164
      ("01", "1000010000111000", "0101110001110110", "0010011111000010"), -- i=1165
      ("10", "1000010000111000", "0101110001110110", "0000010000110000"), -- i=1166
      ("11", "1000010000111000", "0101110001110110", "1101110001111110"), -- i=1167
      ("00", "0100111000000100", "1001101111010110", "1110100111011010"), -- i=1168
      ("01", "0100111000000100", "1001101111010110", "1011001000101110"), -- i=1169
      ("10", "0100111000000100", "1001101111010110", "0000101000000100"), -- i=1170
      ("11", "0100111000000100", "1001101111010110", "1101111111010110"), -- i=1171
      ("00", "1000001111001110", "1010100000001010", "0010101111011000"), -- i=1172
      ("01", "1000001111001110", "1010100000001010", "1101101111000100"), -- i=1173
      ("10", "1000001111001110", "1010100000001010", "1000000000001010"), -- i=1174
      ("11", "1000001111001110", "1010100000001010", "1010101111001110"), -- i=1175
      ("00", "0000101010011100", "1011110100010101", "1100011110110001"), -- i=1176
      ("01", "0000101010011100", "1011110100010101", "0100110110000111"), -- i=1177
      ("10", "0000101010011100", "1011110100010101", "0000100000010100"), -- i=1178
      ("11", "0000101010011100", "1011110100010101", "1011111110011101"), -- i=1179
      ("00", "0010100000110110", "1010000010011010", "1100100011010000"), -- i=1180
      ("01", "0010100000110110", "1010000010011010", "1000011110011100"), -- i=1181
      ("10", "0010100000110110", "1010000010011010", "0010000000010010"), -- i=1182
      ("11", "0010100000110110", "1010000010011010", "1010100010111110"), -- i=1183
      ("00", "1001101000011011", "1011001001001000", "0100110001100011"), -- i=1184
      ("01", "1001101000011011", "1011001001001000", "1110011111010011"), -- i=1185
      ("10", "1001101000011011", "1011001001001000", "1001001000001000"), -- i=1186
      ("11", "1001101000011011", "1011001001001000", "1011101001011011"), -- i=1187
      ("00", "0000010111010101", "1001001111011010", "1001100110101111"), -- i=1188
      ("01", "0000010111010101", "1001001111011010", "0111000111111011"), -- i=1189
      ("10", "0000010111010101", "1001001111011010", "0000000111010000"), -- i=1190
      ("11", "0000010111010101", "1001001111011010", "1001011111011111"), -- i=1191
      ("00", "0101011010100001", "1110001110110100", "0011101001010101"), -- i=1192
      ("01", "0101011010100001", "1110001110110100", "0111001011101101"), -- i=1193
      ("10", "0101011010100001", "1110001110110100", "0100001010100000"), -- i=1194
      ("11", "0101011010100001", "1110001110110100", "1111011110110101"), -- i=1195
      ("00", "1101010110011110", "1110110100010111", "1100001010110101"), -- i=1196
      ("01", "1101010110011110", "1110110100010111", "1110100010000111"), -- i=1197
      ("10", "1101010110011110", "1110110100010111", "1100010100010110"), -- i=1198
      ("11", "1101010110011110", "1110110100010111", "1111110110011111"), -- i=1199
      ("00", "1111001100001110", "0111001100101001", "0110011000110111"), -- i=1200
      ("01", "1111001100001110", "0111001100101001", "0111111111100101"), -- i=1201
      ("10", "1111001100001110", "0111001100101001", "0111001100001000"), -- i=1202
      ("11", "1111001100001110", "0111001100101001", "1111001100101111"), -- i=1203
      ("00", "0000001000100110", "1000110000001111", "1000111000110101"), -- i=1204
      ("01", "0000001000100110", "1000110000001111", "0111011000010111"), -- i=1205
      ("10", "0000001000100110", "1000110000001111", "0000000000000110"), -- i=1206
      ("11", "0000001000100110", "1000110000001111", "1000111000101111"), -- i=1207
      ("00", "1001101011101010", "1000011001010110", "0010000101000000"), -- i=1208
      ("01", "1001101011101010", "1000011001010110", "0001010010010100"), -- i=1209
      ("10", "1001101011101010", "1000011001010110", "1000001001000010"), -- i=1210
      ("11", "1001101011101010", "1000011001010110", "1001111011111110"), -- i=1211
      ("00", "0000011101001101", "1110100000010100", "1110111101100001"), -- i=1212
      ("01", "0000011101001101", "1110100000010100", "0001111100111001"), -- i=1213
      ("10", "0000011101001101", "1110100000010100", "0000000000000100"), -- i=1214
      ("11", "0000011101001101", "1110100000010100", "1110111101011101"), -- i=1215
      ("00", "1000000000110000", "0000101110111111", "1000101111101111"), -- i=1216
      ("01", "1000000000110000", "0000101110111111", "0111010001110001"), -- i=1217
      ("10", "1000000000110000", "0000101110111111", "0000000000110000"), -- i=1218
      ("11", "1000000000110000", "0000101110111111", "1000101110111111"), -- i=1219
      ("00", "0000110010001010", "1011011000010111", "1100001010100001"), -- i=1220
      ("01", "0000110010001010", "1011011000010111", "0101011001110011"), -- i=1221
      ("10", "0000110010001010", "1011011000010111", "0000010000000010"), -- i=1222
      ("11", "0000110010001010", "1011011000010111", "1011111010011111"), -- i=1223
      ("00", "0110011011001100", "0011000110111011", "1001100010000111"), -- i=1224
      ("01", "0110011011001100", "0011000110111011", "0011010100010001"), -- i=1225
      ("10", "0110011011001100", "0011000110111011", "0010000010001000"), -- i=1226
      ("11", "0110011011001100", "0011000110111011", "0111011111111111"), -- i=1227
      ("00", "0100101100110001", "0011001110001101", "0111111010111110"), -- i=1228
      ("01", "0100101100110001", "0011001110001101", "0001011110100100"), -- i=1229
      ("10", "0100101100110001", "0011001110001101", "0000001100000001"), -- i=1230
      ("11", "0100101100110001", "0011001110001101", "0111101110111101"), -- i=1231
      ("00", "0011101010111011", "1010010111101000", "1110000010100011"), -- i=1232
      ("01", "0011101010111011", "1010010111101000", "1001010011010011"), -- i=1233
      ("10", "0011101010111011", "1010010111101000", "0010000010101000"), -- i=1234
      ("11", "0011101010111011", "1010010111101000", "1011111111111011"), -- i=1235
      ("00", "1110001101011010", "1100101101010101", "1010111010101111"), -- i=1236
      ("01", "1110001101011010", "1100101101010101", "0001100000000101"), -- i=1237
      ("10", "1110001101011010", "1100101101010101", "1100001101010000"), -- i=1238
      ("11", "1110001101011010", "1100101101010101", "1110101101011111"), -- i=1239
      ("00", "1010001100000110", "0011101100000000", "1101111000000110"), -- i=1240
      ("01", "1010001100000110", "0011101100000000", "0110100000000110"), -- i=1241
      ("10", "1010001100000110", "0011101100000000", "0010001100000000"), -- i=1242
      ("11", "1010001100000110", "0011101100000000", "1011101100000110"), -- i=1243
      ("00", "1011101100111001", "1000010100001010", "0100000001000011"), -- i=1244
      ("01", "1011101100111001", "1000010100001010", "0011011000101111"), -- i=1245
      ("10", "1011101100111001", "1000010100001010", "1000000100001000"), -- i=1246
      ("11", "1011101100111001", "1000010100001010", "1011111100111011"), -- i=1247
      ("00", "1101000100011100", "1100000111110100", "1001001100010000"), -- i=1248
      ("01", "1101000100011100", "1100000111110100", "0000111100101000"), -- i=1249
      ("10", "1101000100011100", "1100000111110100", "1100000100010100"), -- i=1250
      ("11", "1101000100011100", "1100000111110100", "1101000111111100"), -- i=1251
      ("00", "1110010111111111", "1001001001101101", "0111100001101100"), -- i=1252
      ("01", "1110010111111111", "1001001001101101", "0101001110010010"), -- i=1253
      ("10", "1110010111111111", "1001001001101101", "1000000001101101"), -- i=1254
      ("11", "1110010111111111", "1001001001101101", "1111011111111111"), -- i=1255
      ("00", "1000000100111000", "1011101010110111", "0011101111101111"), -- i=1256
      ("01", "1000000100111000", "1011101010110111", "1100011010000001"), -- i=1257
      ("10", "1000000100111000", "1011101010110111", "1000000000110000"), -- i=1258
      ("11", "1000000100111000", "1011101010110111", "1011101110111111"), -- i=1259
      ("00", "1101100010100101", "0101100111001011", "0011001001110000"), -- i=1260
      ("01", "1101100010100101", "0101100111001011", "0111111011011010"), -- i=1261
      ("10", "1101100010100101", "0101100111001011", "0101100010000001"), -- i=1262
      ("11", "1101100010100101", "0101100111001011", "1101100111101111"), -- i=1263
      ("00", "0011110111011001", "0000000000110010", "0011111000001011"), -- i=1264
      ("01", "0011110111011001", "0000000000110010", "0011110110100111"), -- i=1265
      ("10", "0011110111011001", "0000000000110010", "0000000000010000"), -- i=1266
      ("11", "0011110111011001", "0000000000110010", "0011110111111011"), -- i=1267
      ("00", "0110010000111101", "1000111110001110", "1111001111001011"), -- i=1268
      ("01", "0110010000111101", "1000111110001110", "1101010010101111"), -- i=1269
      ("10", "0110010000111101", "1000111110001110", "0000010000001100"), -- i=1270
      ("11", "0110010000111101", "1000111110001110", "1110111110111111"), -- i=1271
      ("00", "0111110101111000", "1011101000101110", "0011011110100110"), -- i=1272
      ("01", "0111110101111000", "1011101000101110", "1100001101001010"), -- i=1273
      ("10", "0111110101111000", "1011101000101110", "0011100000101000"), -- i=1274
      ("11", "0111110101111000", "1011101000101110", "1111111101111110"), -- i=1275
      ("00", "0000011010010111", "0100110001100101", "0101001011111100"), -- i=1276
      ("01", "0000011010010111", "0100110001100101", "1011101000110010"), -- i=1277
      ("10", "0000011010010111", "0100110001100101", "0000010000000101"), -- i=1278
      ("11", "0000011010010111", "0100110001100101", "0100111011110111"), -- i=1279
      ("00", "0001111100001000", "1010111100111100", "1100111001000100"), -- i=1280
      ("01", "0001111100001000", "1010111100111100", "0110111111001100"), -- i=1281
      ("10", "0001111100001000", "1010111100111100", "0000111100001000"), -- i=1282
      ("11", "0001111100001000", "1010111100111100", "1011111100111100"), -- i=1283
      ("00", "1010001101011111", "1001000010100110", "0011010000000101"), -- i=1284
      ("01", "1010001101011111", "1001000010100110", "0001001010111001"), -- i=1285
      ("10", "1010001101011111", "1001000010100110", "1000000000000110"), -- i=1286
      ("11", "1010001101011111", "1001000010100110", "1011001111111111"), -- i=1287
      ("00", "0001111011101011", "1000011111110001", "1010011011011100"), -- i=1288
      ("01", "0001111011101011", "1000011111110001", "1001011011111010"), -- i=1289
      ("10", "0001111011101011", "1000011111110001", "0000011011100001"), -- i=1290
      ("11", "0001111011101011", "1000011111110001", "1001111111111011"), -- i=1291
      ("00", "0010000100001000", "0101000011011001", "0111000111100001"), -- i=1292
      ("01", "0010000100001000", "0101000011011001", "1101000000101111"), -- i=1293
      ("10", "0010000100001000", "0101000011011001", "0000000000001000"), -- i=1294
      ("11", "0010000100001000", "0101000011011001", "0111000111011001"), -- i=1295
      ("00", "0001101101011011", "1011001111101001", "1100111101000100"), -- i=1296
      ("01", "0001101101011011", "1011001111101001", "0110011101110010"), -- i=1297
      ("10", "0001101101011011", "1011001111101001", "0001001101001001"), -- i=1298
      ("11", "0001101101011011", "1011001111101001", "1011101111111011"), -- i=1299
      ("00", "1011011000100111", "1111101010010101", "1011000010111100"), -- i=1300
      ("01", "1011011000100111", "1111101010010101", "1011101110010010"), -- i=1301
      ("10", "1011011000100111", "1111101010010101", "1011001000000101"), -- i=1302
      ("11", "1011011000100111", "1111101010010101", "1111111010110111"), -- i=1303
      ("00", "0110010010000011", "0110100001111001", "1100110011111100"), -- i=1304
      ("01", "0110010010000011", "0110100001111001", "1111110000001010"), -- i=1305
      ("10", "0110010010000011", "0110100001111001", "0110000000000001"), -- i=1306
      ("11", "0110010010000011", "0110100001111001", "0110110011111011"), -- i=1307
      ("00", "1110110100001000", "0101110000011000", "0100100100100000"), -- i=1308
      ("01", "1110110100001000", "0101110000011000", "1001000011110000"), -- i=1309
      ("10", "1110110100001000", "0101110000011000", "0100110000001000"), -- i=1310
      ("11", "1110110100001000", "0101110000011000", "1111110100011000"), -- i=1311
      ("00", "1110000110111111", "1001111111111011", "1000000110111010"), -- i=1312
      ("01", "1110000110111111", "1001111111111011", "0100000111000100"), -- i=1313
      ("10", "1110000110111111", "1001111111111011", "1000000110111011"), -- i=1314
      ("11", "1110000110111111", "1001111111111011", "1111111111111111"), -- i=1315
      ("00", "1000010010100101", "1111110001001000", "1000000011101101"), -- i=1316
      ("01", "1000010010100101", "1111110001001000", "1000100001011101"), -- i=1317
      ("10", "1000010010100101", "1111110001001000", "1000010000000000"), -- i=1318
      ("11", "1000010010100101", "1111110001001000", "1111110011101101"), -- i=1319
      ("00", "0000101011000010", "0001100000010110", "0010001011011000"), -- i=1320
      ("01", "0000101011000010", "0001100000010110", "1111001010101100"), -- i=1321
      ("10", "0000101011000010", "0001100000010110", "0000100000000010"), -- i=1322
      ("11", "0000101011000010", "0001100000010110", "0001101011010110"), -- i=1323
      ("00", "0101111101010110", "0011110000000000", "1001101101010110"), -- i=1324
      ("01", "0101111101010110", "0011110000000000", "0010001101010110"), -- i=1325
      ("10", "0101111101010110", "0011110000000000", "0001110000000000"), -- i=1326
      ("11", "0101111101010110", "0011110000000000", "0111111101010110"), -- i=1327
      ("00", "1001000010010001", "0000110001111111", "1001110100010000"), -- i=1328
      ("01", "1001000010010001", "0000110001111111", "1000010000010010"), -- i=1329
      ("10", "1001000010010001", "0000110001111111", "0000000000010001"), -- i=1330
      ("11", "1001000010010001", "0000110001111111", "1001110011111111"), -- i=1331
      ("00", "1010000011001111", "0000110011010110", "1010110110100101"), -- i=1332
      ("01", "1010000011001111", "0000110011010110", "1001001111111001"), -- i=1333
      ("10", "1010000011001111", "0000110011010110", "0000000011000110"), -- i=1334
      ("11", "1010000011001111", "0000110011010110", "1010110011011111"), -- i=1335
      ("00", "0001011110011101", "1101001100000101", "1110101010100010"), -- i=1336
      ("01", "0001011110011101", "1101001100000101", "0100010010011000"), -- i=1337
      ("10", "0001011110011101", "1101001100000101", "0001001100000101"), -- i=1338
      ("11", "0001011110011101", "1101001100000101", "1101011110011101"), -- i=1339
      ("00", "1111011001001010", "1010010011001011", "1001101100010101"), -- i=1340
      ("01", "1111011001001010", "1010010011001011", "0101000101111111"), -- i=1341
      ("10", "1111011001001010", "1010010011001011", "1010010001001010"), -- i=1342
      ("11", "1111011001001010", "1010010011001011", "1111011011001011"), -- i=1343
      ("00", "1001000101100101", "1000110011100101", "0001111001001010"), -- i=1344
      ("01", "1001000101100101", "1000110011100101", "0000010010000000"), -- i=1345
      ("10", "1001000101100101", "1000110011100101", "1000000001100101"), -- i=1346
      ("11", "1001000101100101", "1000110011100101", "1001110111100101"), -- i=1347
      ("00", "1100010011111001", "0101100110000010", "0001111001111011"), -- i=1348
      ("01", "1100010011111001", "0101100110000010", "0110101101110111"), -- i=1349
      ("10", "1100010011111001", "0101100110000010", "0100000010000000"), -- i=1350
      ("11", "1100010011111001", "0101100110000010", "1101110111111011"), -- i=1351
      ("00", "0101100101101010", "1101100011000010", "0011001000101100"), -- i=1352
      ("01", "0101100101101010", "1101100011000010", "1000000010101000"), -- i=1353
      ("10", "0101100101101010", "1101100011000010", "0101100001000010"), -- i=1354
      ("11", "0101100101101010", "1101100011000010", "1101100111101010"), -- i=1355
      ("00", "1010010000010101", "1011100011110010", "0101110100000111"), -- i=1356
      ("01", "1010010000010101", "1011100011110010", "1110101100100011"), -- i=1357
      ("10", "1010010000010101", "1011100011110010", "1010000000010000"), -- i=1358
      ("11", "1010010000010101", "1011100011110010", "1011110011110111"), -- i=1359
      ("00", "0011011001100010", "1100111111000001", "0000011000100011"), -- i=1360
      ("01", "0011011001100010", "1100111111000001", "0110011010100001"), -- i=1361
      ("10", "0011011001100010", "1100111111000001", "0000011001000000"), -- i=1362
      ("11", "0011011001100010", "1100111111000001", "1111111111100011"), -- i=1363
      ("00", "0001100100100010", "0000100010111100", "0010000111011110"), -- i=1364
      ("01", "0001100100100010", "0000100010111100", "0001000001100110"), -- i=1365
      ("10", "0001100100100010", "0000100010111100", "0000100000100000"), -- i=1366
      ("11", "0001100100100010", "0000100010111100", "0001100110111110"), -- i=1367
      ("00", "1100010111101010", "1001111110001001", "0110010101110011"), -- i=1368
      ("01", "1100010111101010", "1001111110001001", "0010011001100001"), -- i=1369
      ("10", "1100010111101010", "1001111110001001", "1000010110001000"), -- i=1370
      ("11", "1100010111101010", "1001111110001001", "1101111111101011"), -- i=1371
      ("00", "0000011001010010", "1001000010000110", "1001011011011000"), -- i=1372
      ("01", "0000011001010010", "1001000010000110", "0111010111001100"), -- i=1373
      ("10", "0000011001010010", "1001000010000110", "0000000000000010"), -- i=1374
      ("11", "0000011001010010", "1001000010000110", "1001011011010110"), -- i=1375
      ("00", "1010011000110011", "1100001001001110", "0110100010000001"), -- i=1376
      ("01", "1010011000110011", "1100001001001110", "1110001111100101"), -- i=1377
      ("10", "1010011000110011", "1100001001001110", "1000001000000010"), -- i=1378
      ("11", "1010011000110011", "1100001001001110", "1110011001111111"), -- i=1379
      ("00", "1001110000001001", "0111011100010011", "0001001100011100"), -- i=1380
      ("01", "1001110000001001", "0111011100010011", "0010010011110110"), -- i=1381
      ("10", "1001110000001001", "0111011100010011", "0001010000000001"), -- i=1382
      ("11", "1001110000001001", "0111011100010011", "1111111100011011"), -- i=1383
      ("00", "1110011001011101", "0010110100001100", "0001001101101001"), -- i=1384
      ("01", "1110011001011101", "0010110100001100", "1011100101010001"), -- i=1385
      ("10", "1110011001011101", "0010110100001100", "0010010000001100"), -- i=1386
      ("11", "1110011001011101", "0010110100001100", "1110111101011101"), -- i=1387
      ("00", "1110011111101111", "1000010011110111", "0110110011100110"), -- i=1388
      ("01", "1110011111101111", "1000010011110111", "0110001011111000"), -- i=1389
      ("10", "1110011111101111", "1000010011110111", "1000010011100111"), -- i=1390
      ("11", "1110011111101111", "1000010011110111", "1110011111111111"), -- i=1391
      ("00", "1110001110000111", "1100101110011100", "1010111100100011"), -- i=1392
      ("01", "1110001110000111", "1100101110011100", "0001011111101011"), -- i=1393
      ("10", "1110001110000111", "1100101110011100", "1100001110000100"), -- i=1394
      ("11", "1110001110000111", "1100101110011100", "1110101110011111"), -- i=1395
      ("00", "0100110100100011", "1101001100010111", "0010000000111010"), -- i=1396
      ("01", "0100110100100011", "1101001100010111", "0111101000001100"), -- i=1397
      ("10", "0100110100100011", "1101001100010111", "0100000100000011"), -- i=1398
      ("11", "0100110100100011", "1101001100010111", "1101111100110111"), -- i=1399
      ("00", "1011110110110110", "0100100101011100", "0000011100010010"), -- i=1400
      ("01", "1011110110110110", "0100100101011100", "0111010001011010"), -- i=1401
      ("10", "1011110110110110", "0100100101011100", "0000100100010100"), -- i=1402
      ("11", "1011110110110110", "0100100101011100", "1111110111111110"), -- i=1403
      ("00", "0100101001100110", "0100011001011001", "1001000010111111"), -- i=1404
      ("01", "0100101001100110", "0100011001011001", "0000010000001101"), -- i=1405
      ("10", "0100101001100110", "0100011001011001", "0100001001000000"), -- i=1406
      ("11", "0100101001100110", "0100011001011001", "0100111001111111"), -- i=1407
      ("00", "1111110100101111", "0111010001110100", "0111000110100011"), -- i=1408
      ("01", "1111110100101111", "0111010001110100", "1000100010111011"), -- i=1409
      ("10", "1111110100101111", "0111010001110100", "0111010000100100"), -- i=1410
      ("11", "1111110100101111", "0111010001110100", "1111110101111111"), -- i=1411
      ("00", "1111010001100000", "1011110100110111", "1011000110010111"), -- i=1412
      ("01", "1111010001100000", "1011110100110111", "0011011100101001"), -- i=1413
      ("10", "1111010001100000", "1011110100110111", "1011010000100000"), -- i=1414
      ("11", "1111010001100000", "1011110100110111", "1111110101110111"), -- i=1415
      ("00", "1101010111011001", "1000000100001011", "0101011011100100"), -- i=1416
      ("01", "1101010111011001", "1000000100001011", "0101010011001110"), -- i=1417
      ("10", "1101010111011001", "1000000100001011", "1000000100001001"), -- i=1418
      ("11", "1101010111011001", "1000000100001011", "1101010111011011"), -- i=1419
      ("00", "0111001101001101", "1111111100010011", "0111001001100000"), -- i=1420
      ("01", "0111001101001101", "1111111100010011", "0111010000111010"), -- i=1421
      ("10", "0111001101001101", "1111111100010011", "0111001100000001"), -- i=1422
      ("11", "0111001101001101", "1111111100010011", "1111111101011111"), -- i=1423
      ("00", "1011001111000011", "0001000011101111", "1100010010110010"), -- i=1424
      ("01", "1011001111000011", "0001000011101111", "1010001011010100"), -- i=1425
      ("10", "1011001111000011", "0001000011101111", "0001000011000011"), -- i=1426
      ("11", "1011001111000011", "0001000011101111", "1011001111101111"), -- i=1427
      ("00", "1010010011000000", "1101000010001001", "0111010101001001"), -- i=1428
      ("01", "1010010011000000", "1101000010001001", "1101010000110111"), -- i=1429
      ("10", "1010010011000000", "1101000010001001", "1000000010000000"), -- i=1430
      ("11", "1010010011000000", "1101000010001001", "1111010011001001"), -- i=1431
      ("00", "0110000011110000", "0010101101111010", "1000110001101010"), -- i=1432
      ("01", "0110000011110000", "0010101101111010", "0011010101110110"), -- i=1433
      ("10", "0110000011110000", "0010101101111010", "0010000001110000"), -- i=1434
      ("11", "0110000011110000", "0010101101111010", "0110101111111010"), -- i=1435
      ("00", "1011101100111000", "0000101100001001", "1100011001000001"), -- i=1436
      ("01", "1011101100111000", "0000101100001001", "1011000000101111"), -- i=1437
      ("10", "1011101100111000", "0000101100001001", "0000101100001000"), -- i=1438
      ("11", "1011101100111000", "0000101100001001", "1011101100111001"), -- i=1439
      ("00", "0010000111101000", "0100000011000101", "0110001010101101"), -- i=1440
      ("01", "0010000111101000", "0100000011000101", "1110000100100011"), -- i=1441
      ("10", "0010000111101000", "0100000011000101", "0000000011000000"), -- i=1442
      ("11", "0010000111101000", "0100000011000101", "0110000111101101"), -- i=1443
      ("00", "0101011011000100", "0011100110001111", "1001000001010011"), -- i=1444
      ("01", "0101011011000100", "0011100110001111", "0001110100110101"), -- i=1445
      ("10", "0101011011000100", "0011100110001111", "0001000010000100"), -- i=1446
      ("11", "0101011011000100", "0011100110001111", "0111111111001111"), -- i=1447
      ("00", "1001101111011000", "1110101001100100", "1000011000111100"), -- i=1448
      ("01", "1001101111011000", "1110101001100100", "1011000101110100"), -- i=1449
      ("10", "1001101111011000", "1110101001100100", "1000101001000000"), -- i=1450
      ("11", "1001101111011000", "1110101001100100", "1111101111111100"), -- i=1451
      ("00", "0001101011110000", "0000011100110101", "0010001000100101"), -- i=1452
      ("01", "0001101011110000", "0000011100110101", "0001001110111011"), -- i=1453
      ("10", "0001101011110000", "0000011100110101", "0000001000110000"), -- i=1454
      ("11", "0001101011110000", "0000011100110101", "0001111111110101"), -- i=1455
      ("00", "0011010000100000", "0101101101001100", "1000111101101100"), -- i=1456
      ("01", "0011010000100000", "0101101101001100", "1101100011010100"), -- i=1457
      ("10", "0011010000100000", "0101101101001100", "0001000000000000"), -- i=1458
      ("11", "0011010000100000", "0101101101001100", "0111111101101100"), -- i=1459
      ("00", "0011011110101101", "1011111111101100", "1111011110011001"), -- i=1460
      ("01", "0011011110101101", "1011111111101100", "0111011111000001"), -- i=1461
      ("10", "0011011110101101", "1011111111101100", "0011011110101100"), -- i=1462
      ("11", "0011011110101101", "1011111111101100", "1011111111101101"), -- i=1463
      ("00", "1101111010011111", "0101011110010100", "0011011000110011"), -- i=1464
      ("01", "1101111010011111", "0101011110010100", "1000011100001011"), -- i=1465
      ("10", "1101111010011111", "0101011110010100", "0101011010010100"), -- i=1466
      ("11", "1101111010011111", "0101011110010100", "1101111110011111"), -- i=1467
      ("00", "1011001111111111", "0011111010110111", "1111001010110110"), -- i=1468
      ("01", "1011001111111111", "0011111010110111", "0111010101001000"), -- i=1469
      ("10", "1011001111111111", "0011111010110111", "0011001010110111"), -- i=1470
      ("11", "1011001111111111", "0011111010110111", "1011111111111111"), -- i=1471
      ("00", "1111110100110001", "0001110000101101", "0001100101011110"), -- i=1472
      ("01", "1111110100110001", "0001110000101101", "1110000100000100"), -- i=1473
      ("10", "1111110100110001", "0001110000101101", "0001110000100001"), -- i=1474
      ("11", "1111110100110001", "0001110000101101", "1111110100111101"), -- i=1475
      ("00", "1000101010010000", "1110100000001101", "0111001010011101"), -- i=1476
      ("01", "1000101010010000", "1110100000001101", "1010001010000011"), -- i=1477
      ("10", "1000101010010000", "1110100000001101", "1000100000000000"), -- i=1478
      ("11", "1000101010010000", "1110100000001101", "1110101010011101"), -- i=1479
      ("00", "0000100000010010", "1101010111010101", "1101110111100111"), -- i=1480
      ("01", "0000100000010010", "1101010111010101", "0011001000111101"), -- i=1481
      ("10", "0000100000010010", "1101010111010101", "0000000000010000"), -- i=1482
      ("11", "0000100000010010", "1101010111010101", "1101110111010111"), -- i=1483
      ("00", "1101000110001011", "1011101001011011", "1000101111100110"), -- i=1484
      ("01", "1101000110001011", "1011101001011011", "0001011100110000"), -- i=1485
      ("10", "1101000110001011", "1011101001011011", "1001000000001011"), -- i=1486
      ("11", "1101000110001011", "1011101001011011", "1111101111011011"), -- i=1487
      ("00", "0011010000100110", "0010010111001011", "0101100111110001"), -- i=1488
      ("01", "0011010000100110", "0010010111001011", "0000111001011011"), -- i=1489
      ("10", "0011010000100110", "0010010111001011", "0010010000000010"), -- i=1490
      ("11", "0011010000100110", "0010010111001011", "0011010111101111"), -- i=1491
      ("00", "0011100001000000", "0001000111000011", "0100101000000011"), -- i=1492
      ("01", "0011100001000000", "0001000111000011", "0010011001111101"), -- i=1493
      ("10", "0011100001000000", "0001000111000011", "0001000001000000"), -- i=1494
      ("11", "0011100001000000", "0001000111000011", "0011100111000011"), -- i=1495
      ("00", "0011000101100101", "1011101000010101", "1110101101111010"), -- i=1496
      ("01", "0011000101100101", "1011101000010101", "0111011101010000"), -- i=1497
      ("10", "0011000101100101", "1011101000010101", "0011000000000101"), -- i=1498
      ("11", "0011000101100101", "1011101000010101", "1011101101110101"), -- i=1499
      ("00", "0001111010001110", "0111011110001011", "1001011000011001"), -- i=1500
      ("01", "0001111010001110", "0111011110001011", "1010011100000011"), -- i=1501
      ("10", "0001111010001110", "0111011110001011", "0001011010001010"), -- i=1502
      ("11", "0001111010001110", "0111011110001011", "0111111110001111"), -- i=1503
      ("00", "0110100011011000", "0010111001011110", "1001011100110110"), -- i=1504
      ("01", "0110100011011000", "0010111001011110", "0011101001111010"), -- i=1505
      ("10", "0110100011011000", "0010111001011110", "0010100001011000"), -- i=1506
      ("11", "0110100011011000", "0010111001011110", "0110111011011110"), -- i=1507
      ("00", "0110101100001011", "1011100011011011", "0010001111100110"), -- i=1508
      ("01", "0110101100001011", "1011100011011011", "1011001000110000"), -- i=1509
      ("10", "0110101100001011", "1011100011011011", "0010100000001011"), -- i=1510
      ("11", "0110101100001011", "1011100011011011", "1111101111011011"), -- i=1511
      ("00", "1101011011101101", "0100000110111001", "0001100010100110"), -- i=1512
      ("01", "1101011011101101", "0100000110111001", "1001010100110100"), -- i=1513
      ("10", "1101011011101101", "0100000110111001", "0100000010101001"), -- i=1514
      ("11", "1101011011101101", "0100000110111001", "1101011111111101"), -- i=1515
      ("00", "0000111001011011", "1000101111000001", "1001101000011100"), -- i=1516
      ("01", "0000111001011011", "1000101111000001", "1000001010011010"), -- i=1517
      ("10", "0000111001011011", "1000101111000001", "0000101001000001"), -- i=1518
      ("11", "0000111001011011", "1000101111000001", "1000111111011011"), -- i=1519
      ("00", "1011110000010111", "1110110011001010", "1010100011100001"), -- i=1520
      ("01", "1011110000010111", "1110110011001010", "1100111101001101"), -- i=1521
      ("10", "1011110000010111", "1110110011001010", "1010110000000010"), -- i=1522
      ("11", "1011110000010111", "1110110011001010", "1111110011011111"), -- i=1523
      ("00", "1101001101001001", "0011110010011100", "0000111111100101"), -- i=1524
      ("01", "1101001101001001", "0011110010011100", "1001011010101101"), -- i=1525
      ("10", "1101001101001001", "0011110010011100", "0001000000001000"), -- i=1526
      ("11", "1101001101001001", "0011110010011100", "1111111111011101"), -- i=1527
      ("00", "1110001011101111", "0000101100101101", "1110111000011100"), -- i=1528
      ("01", "1110001011101111", "0000101100101101", "1101011111000010"), -- i=1529
      ("10", "1110001011101111", "0000101100101101", "0000001000101101"), -- i=1530
      ("11", "1110001011101111", "0000101100101101", "1110101111101111"), -- i=1531
      ("00", "1011010001110110", "0011100101011111", "1110110111010101"), -- i=1532
      ("01", "1011010001110110", "0011100101011111", "0111101100010111"), -- i=1533
      ("10", "1011010001110110", "0011100101011111", "0011000001010110"), -- i=1534
      ("11", "1011010001110110", "0011100101011111", "1011110101111111"), -- i=1535
      ("00", "0010100001011111", "0001101000011011", "0100001001111010"), -- i=1536
      ("01", "0010100001011111", "0001101000011011", "0000111001000100"), -- i=1537
      ("10", "0010100001011111", "0001101000011011", "0000100000011011"), -- i=1538
      ("11", "0010100001011111", "0001101000011011", "0011101001011111"), -- i=1539
      ("00", "0111000111000011", "1101001101001000", "0100010100001011"), -- i=1540
      ("01", "0111000111000011", "1101001101001000", "1001111001111011"), -- i=1541
      ("10", "0111000111000011", "1101001101001000", "0101000101000000"), -- i=1542
      ("11", "0111000111000011", "1101001101001000", "1111001111001011"), -- i=1543
      ("00", "0100011101111111", "0000010110011010", "0100110100011001"), -- i=1544
      ("01", "0100011101111111", "0000010110011010", "0100000111100101"), -- i=1545
      ("10", "0100011101111111", "0000010110011010", "0000010100011010"), -- i=1546
      ("11", "0100011101111111", "0000010110011010", "0100011111111111"), -- i=1547
      ("00", "1000100011000110", "0011101100001001", "1100001111001111"), -- i=1548
      ("01", "1000100011000110", "0011101100001001", "0100110110111101"), -- i=1549
      ("10", "1000100011000110", "0011101100001001", "0000100000000000"), -- i=1550
      ("11", "1000100011000110", "0011101100001001", "1011101111001111"), -- i=1551
      ("00", "1010100000101000", "0001110011000010", "1100010011101010"), -- i=1552
      ("01", "1010100000101000", "0001110011000010", "1000101101100110"), -- i=1553
      ("10", "1010100000101000", "0001110011000010", "0000100000000000"), -- i=1554
      ("11", "1010100000101000", "0001110011000010", "1011110011101010"), -- i=1555
      ("00", "0000010011101100", "1000111010000000", "1001001101101100"), -- i=1556
      ("01", "0000010011101100", "1000111010000000", "0111011001101100"), -- i=1557
      ("10", "0000010011101100", "1000111010000000", "0000010010000000"), -- i=1558
      ("11", "0000010011101100", "1000111010000000", "1000111011101100"), -- i=1559
      ("00", "0001010001111000", "0000110011011111", "0010000101010111"), -- i=1560
      ("01", "0001010001111000", "0000110011011111", "0000011110011001"), -- i=1561
      ("10", "0001010001111000", "0000110011011111", "0000010001011000"), -- i=1562
      ("11", "0001010001111000", "0000110011011111", "0001110011111111"), -- i=1563
      ("00", "1101010100011000", "1100101001101000", "1001111110000000"), -- i=1564
      ("01", "1101010100011000", "1100101001101000", "0000101010110000"), -- i=1565
      ("10", "1101010100011000", "1100101001101000", "1100000000001000"), -- i=1566
      ("11", "1101010100011000", "1100101001101000", "1101111101111000"), -- i=1567
      ("00", "1100011010111101", "0011001010000000", "1111100100111101"), -- i=1568
      ("01", "1100011010111101", "0011001010000000", "1001010000111101"), -- i=1569
      ("10", "1100011010111101", "0011001010000000", "0000001010000000"), -- i=1570
      ("11", "1100011010111101", "0011001010000000", "1111011010111101"), -- i=1571
      ("00", "0111010111101010", "1001010110101111", "0000101110011001"), -- i=1572
      ("01", "0111010111101010", "1001010110101111", "1110000000111011"), -- i=1573
      ("10", "0111010111101010", "1001010110101111", "0001010110101010"), -- i=1574
      ("11", "0111010111101010", "1001010110101111", "1111010111101111"), -- i=1575
      ("00", "0011011010000100", "1010011010110100", "1101110100111000"), -- i=1576
      ("01", "0011011010000100", "1010011010110100", "1000111111010000"), -- i=1577
      ("10", "0011011010000100", "1010011010110100", "0010011010000100"), -- i=1578
      ("11", "0011011010000100", "1010011010110100", "1011011010110100"), -- i=1579
      ("00", "1100100011110010", "0010011101100110", "1111000001011000"), -- i=1580
      ("01", "1100100011110010", "0010011101100110", "1010000110001100"), -- i=1581
      ("10", "1100100011110010", "0010011101100110", "0000000001100010"), -- i=1582
      ("11", "1100100011110010", "0010011101100110", "1110111111110110"), -- i=1583
      ("00", "0110100010111011", "0010111000001000", "1001011011000011"), -- i=1584
      ("01", "0110100010111011", "0010111000001000", "0011101010110011"), -- i=1585
      ("10", "0110100010111011", "0010111000001000", "0010100000001000"), -- i=1586
      ("11", "0110100010111011", "0010111000001000", "0110111010111011"), -- i=1587
      ("00", "1110001001111011", "1111101101011001", "1101110111010100"), -- i=1588
      ("01", "1110001001111011", "1111101101011001", "1110011100100010"), -- i=1589
      ("10", "1110001001111011", "1111101101011001", "1110001001011001"), -- i=1590
      ("11", "1110001001111011", "1111101101011001", "1111101101111011"), -- i=1591
      ("00", "0100110000111011", "1001011000000110", "1110001001000001"), -- i=1592
      ("01", "0100110000111011", "1001011000000110", "1011011000110101"), -- i=1593
      ("10", "0100110000111011", "1001011000000110", "0000010000000010"), -- i=1594
      ("11", "0100110000111011", "1001011000000110", "1101111000111111"), -- i=1595
      ("00", "0111000011000010", "1010010011011111", "0001010110100001"), -- i=1596
      ("01", "0111000011000010", "1010010011011111", "1100101111100011"), -- i=1597
      ("10", "0111000011000010", "1010010011011111", "0010000011000010"), -- i=1598
      ("11", "0111000011000010", "1010010011011111", "1111010011011111"), -- i=1599
      ("00", "1101100100010000", "0001110101001111", "1111011001011111"), -- i=1600
      ("01", "1101100100010000", "0001110101001111", "1011101111000001"), -- i=1601
      ("10", "1101100100010000", "0001110101001111", "0001100100000000"), -- i=1602
      ("11", "1101100100010000", "0001110101001111", "1101110101011111"), -- i=1603
      ("00", "0010000010101010", "1101001001100110", "1111001100010000"), -- i=1604
      ("01", "0010000010101010", "1101001001100110", "0100111001000100"), -- i=1605
      ("10", "0010000010101010", "1101001001100110", "0000000000100010"), -- i=1606
      ("11", "0010000010101010", "1101001001100110", "1111001011101110"), -- i=1607
      ("00", "0011111001010111", "0011100110000100", "0111011111011011"), -- i=1608
      ("01", "0011111001010111", "0011100110000100", "0000010011010011"), -- i=1609
      ("10", "0011111001010111", "0011100110000100", "0011100000000100"), -- i=1610
      ("11", "0011111001010111", "0011100110000100", "0011111111010111"), -- i=1611
      ("00", "0000110101011011", "0111111111000011", "1000110100011110"), -- i=1612
      ("01", "0000110101011011", "0111111111000011", "1000110110011000"), -- i=1613
      ("10", "0000110101011011", "0111111111000011", "0000110101000011"), -- i=1614
      ("11", "0000110101011011", "0111111111000011", "0111111111011011"), -- i=1615
      ("00", "0110011110011011", "0110110110011011", "1101010100110110"), -- i=1616
      ("01", "0110011110011011", "0110110110011011", "1111101000000000"), -- i=1617
      ("10", "0110011110011011", "0110110110011011", "0110010110011011"), -- i=1618
      ("11", "0110011110011011", "0110110110011011", "0110111110011011"), -- i=1619
      ("00", "1101100101010011", "0110100001011111", "0100000110110010"), -- i=1620
      ("01", "1101100101010011", "0110100001011111", "0111000011110100"), -- i=1621
      ("10", "1101100101010011", "0110100001011111", "0100100001010011"), -- i=1622
      ("11", "1101100101010011", "0110100001011111", "1111100101011111"), -- i=1623
      ("00", "1000011111110101", "1110101001100001", "0111001001010110"), -- i=1624
      ("01", "1000011111110101", "1110101001100001", "1001110110010100"), -- i=1625
      ("10", "1000011111110101", "1110101001100001", "1000001001100001"), -- i=1626
      ("11", "1000011111110101", "1110101001100001", "1110111111110101"), -- i=1627
      ("00", "1000100011001010", "0000010110101110", "1000111001111000"), -- i=1628
      ("01", "1000100011001010", "0000010110101110", "1000001100011100"), -- i=1629
      ("10", "1000100011001010", "0000010110101110", "0000000010001010"), -- i=1630
      ("11", "1000100011001010", "0000010110101110", "1000110111101110"), -- i=1631
      ("00", "0010011001011011", "0110001000111000", "1000100010010011"), -- i=1632
      ("01", "0010011001011011", "0110001000111000", "1100010000100011"), -- i=1633
      ("10", "0010011001011011", "0110001000111000", "0010001000011000"), -- i=1634
      ("11", "0010011001011011", "0110001000111000", "0110011001111011"), -- i=1635
      ("00", "1001011010000110", "1100100110100001", "0110000000100111"), -- i=1636
      ("01", "1001011010000110", "1100100110100001", "1100110011100101"), -- i=1637
      ("10", "1001011010000110", "1100100110100001", "1000000010000000"), -- i=1638
      ("11", "1001011010000110", "1100100110100001", "1101111110100111"), -- i=1639
      ("00", "0101101111110001", "1101000001001110", "0010110000111111"), -- i=1640
      ("01", "0101101111110001", "1101000001001110", "1000101110100011"), -- i=1641
      ("10", "0101101111110001", "1101000001001110", "0101000001000000"), -- i=1642
      ("11", "0101101111110001", "1101000001001110", "1101101111111111"), -- i=1643
      ("00", "0000010101110111", "1100111111110010", "1101010101101001"), -- i=1644
      ("01", "0000010101110111", "1100111111110010", "0011010110000101"), -- i=1645
      ("10", "0000010101110111", "1100111111110010", "0000010101110010"), -- i=1646
      ("11", "0000010101110111", "1100111111110010", "1100111111110111"), -- i=1647
      ("00", "1001001000110011", "1111001011101110", "1000010100100001"), -- i=1648
      ("01", "1001001000110011", "1111001011101110", "1001111101000101"), -- i=1649
      ("10", "1001001000110011", "1111001011101110", "1001001000100010"), -- i=1650
      ("11", "1001001000110011", "1111001011101110", "1111001011111111"), -- i=1651
      ("00", "0110001010110010", "1111010010000000", "0101011100110010"), -- i=1652
      ("01", "0110001010110010", "1111010010000000", "0110111000110010"), -- i=1653
      ("10", "0110001010110010", "1111010010000000", "0110000010000000"), -- i=1654
      ("11", "0110001010110010", "1111010010000000", "1111011010110010"), -- i=1655
      ("00", "0001010001010110", "1101111110011110", "1111001111110100"), -- i=1656
      ("01", "0001010001010110", "1101111110011110", "0011010010111000"), -- i=1657
      ("10", "0001010001010110", "1101111110011110", "0001010000010110"), -- i=1658
      ("11", "0001010001010110", "1101111110011110", "1101111111011110"), -- i=1659
      ("00", "1100010010100111", "0001100000011000", "1101110010111111"), -- i=1660
      ("01", "1100010010100111", "0001100000011000", "1010110010001111"), -- i=1661
      ("10", "1100010010100111", "0001100000011000", "0000000000000000"), -- i=1662
      ("11", "1100010010100111", "0001100000011000", "1101110010111111"), -- i=1663
      ("00", "0011010001000000", "0110011100100010", "1001101101100010"), -- i=1664
      ("01", "0011010001000000", "0110011100100010", "1100110100011110"), -- i=1665
      ("10", "0011010001000000", "0110011100100010", "0010010000000000"), -- i=1666
      ("11", "0011010001000000", "0110011100100010", "0111011101100010"), -- i=1667
      ("00", "1101010110101111", "0110000001100010", "0011011000010001"), -- i=1668
      ("01", "1101010110101111", "0110000001100010", "0111010101001101"), -- i=1669
      ("10", "1101010110101111", "0110000001100010", "0100000000100010"), -- i=1670
      ("11", "1101010110101111", "0110000001100010", "1111010111101111"), -- i=1671
      ("00", "1001100011011110", "1111011010101010", "1000111110001000"), -- i=1672
      ("01", "1001100011011110", "1111011010101010", "1010001000110100"), -- i=1673
      ("10", "1001100011011110", "1111011010101010", "1001000010001010"), -- i=1674
      ("11", "1001100011011110", "1111011010101010", "1111111011111110"), -- i=1675
      ("00", "1110000101000110", "0110101011010001", "0100110000010111"), -- i=1676
      ("01", "1110000101000110", "0110101011010001", "0111011001110101"), -- i=1677
      ("10", "1110000101000110", "0110101011010001", "0110000001000000"), -- i=1678
      ("11", "1110000101000110", "0110101011010001", "1110101111010111"), -- i=1679
      ("00", "1000100011001001", "0100001010110001", "1100101101111010"), -- i=1680
      ("01", "1000100011001001", "0100001010110001", "0100011000011000"), -- i=1681
      ("10", "1000100011001001", "0100001010110001", "0000000010000001"), -- i=1682
      ("11", "1000100011001001", "0100001010110001", "1100101011111001"), -- i=1683
      ("00", "1010110010010010", "1011110111001011", "0110101001011101"), -- i=1684
      ("01", "1010110010010010", "1011110111001011", "1110111011000111"), -- i=1685
      ("10", "1010110010010010", "1011110111001011", "1010110010000010"), -- i=1686
      ("11", "1010110010010010", "1011110111001011", "1011110111011011"), -- i=1687
      ("00", "1010100110000101", "0100111101100001", "1111100011100110"), -- i=1688
      ("01", "1010100110000101", "0100111101100001", "0101101000100100"), -- i=1689
      ("10", "1010100110000101", "0100111101100001", "0000100100000001"), -- i=1690
      ("11", "1010100110000101", "0100111101100001", "1110111111100101"), -- i=1691
      ("00", "1001110000001011", "0011111001100010", "1101101001101101"), -- i=1692
      ("01", "1001110000001011", "0011111001100010", "0101110110101001"), -- i=1693
      ("10", "1001110000001011", "0011111001100010", "0001110000000010"), -- i=1694
      ("11", "1001110000001011", "0011111001100010", "1011111001101011"), -- i=1695
      ("00", "1011100010111001", "0101100101111010", "0001001000110011"), -- i=1696
      ("01", "1011100010111001", "0101100101111010", "0101111100111111"), -- i=1697
      ("10", "1011100010111001", "0101100101111010", "0001100000111000"), -- i=1698
      ("11", "1011100010111001", "0101100101111010", "1111100111111011"), -- i=1699
      ("00", "0100100101011111", "0001010001011111", "0101110110111110"), -- i=1700
      ("01", "0100100101011111", "0001010001011111", "0011010100000000"), -- i=1701
      ("10", "0100100101011111", "0001010001011111", "0000000001011111"), -- i=1702
      ("11", "0100100101011111", "0001010001011111", "0101110101011111"), -- i=1703
      ("00", "0011101000111000", "1011101000001110", "1111010001000110"), -- i=1704
      ("01", "0011101000111000", "1011101000001110", "1000000000101010"), -- i=1705
      ("10", "0011101000111000", "1011101000001110", "0011101000001000"), -- i=1706
      ("11", "0011101000111000", "1011101000001110", "1011101000111110"), -- i=1707
      ("00", "0011010111110001", "0011000101111000", "0110011101101001"), -- i=1708
      ("01", "0011010111110001", "0011000101111000", "0000010001111001"), -- i=1709
      ("10", "0011010111110001", "0011000101111000", "0011000101110000"), -- i=1710
      ("11", "0011010111110001", "0011000101111000", "0011010111111001"), -- i=1711
      ("00", "1111001010111001", "0001111010011101", "0001000101010110"), -- i=1712
      ("01", "1111001010111001", "0001111010011101", "1101010000011100"), -- i=1713
      ("10", "1111001010111001", "0001111010011101", "0001001010011001"), -- i=1714
      ("11", "1111001010111001", "0001111010011101", "1111111010111101"), -- i=1715
      ("00", "1011011110000101", "1010001111011001", "0101101101011110"), -- i=1716
      ("01", "1011011110000101", "1010001111011001", "0001001110101100"), -- i=1717
      ("10", "1011011110000101", "1010001111011001", "1010001110000001"), -- i=1718
      ("11", "1011011110000101", "1010001111011001", "1011011111011101"), -- i=1719
      ("00", "0100110010010000", "0101011001010010", "1010001011100010"), -- i=1720
      ("01", "0100110010010000", "0101011001010010", "1111011000111110"), -- i=1721
      ("10", "0100110010010000", "0101011001010010", "0100010000010000"), -- i=1722
      ("11", "0100110010010000", "0101011001010010", "0101111011010010"), -- i=1723
      ("00", "1001010111111101", "1111011101111110", "1000110101111011"), -- i=1724
      ("01", "1001010111111101", "1111011101111110", "1001111001111111"), -- i=1725
      ("10", "1001010111111101", "1111011101111110", "1001010101111100"), -- i=1726
      ("11", "1001010111111101", "1111011101111110", "1111011111111111"), -- i=1727
      ("00", "0111000011010010", "1000010001110101", "1111010101000111"), -- i=1728
      ("01", "0111000011010010", "1000010001110101", "1110110001011101"), -- i=1729
      ("10", "0111000011010010", "1000010001110101", "0000000001010000"), -- i=1730
      ("11", "0111000011010010", "1000010001110101", "1111010011110111"), -- i=1731
      ("00", "0001001000110101", "0010110011110000", "0011111100100101"), -- i=1732
      ("01", "0001001000110101", "0010110011110000", "1110010101000101"), -- i=1733
      ("10", "0001001000110101", "0010110011110000", "0000000000110000"), -- i=1734
      ("11", "0001001000110101", "0010110011110000", "0011111011110101"), -- i=1735
      ("00", "1111010010100011", "1011111101010101", "1011001111111000"), -- i=1736
      ("01", "1111010010100011", "1011111101010101", "0011010101001110"), -- i=1737
      ("10", "1111010010100011", "1011111101010101", "1011010000000001"), -- i=1738
      ("11", "1111010010100011", "1011111101010101", "1111111111110111"), -- i=1739
      ("00", "0011011101100011", "0011011101011111", "0110111011000010"), -- i=1740
      ("01", "0011011101100011", "0011011101011111", "0000000000000100"), -- i=1741
      ("10", "0011011101100011", "0011011101011111", "0011011101000011"), -- i=1742
      ("11", "0011011101100011", "0011011101011111", "0011011101111111"), -- i=1743
      ("00", "0111011110101101", "0000001000111010", "0111100111100111"), -- i=1744
      ("01", "0111011110101101", "0000001000111010", "0111010101110011"), -- i=1745
      ("10", "0111011110101101", "0000001000111010", "0000001000101000"), -- i=1746
      ("11", "0111011110101101", "0000001000111010", "0111011110111111"), -- i=1747
      ("00", "0110100110001100", "1000011100111001", "1111000011000101"), -- i=1748
      ("01", "0110100110001100", "1000011100111001", "1110001001010011"), -- i=1749
      ("10", "0110100110001100", "1000011100111001", "0000000100001000"), -- i=1750
      ("11", "0110100110001100", "1000011100111001", "1110111110111101"), -- i=1751
      ("00", "0111010111101110", "1110000000100100", "0101011000010010"), -- i=1752
      ("01", "0111010111101110", "1110000000100100", "1001010111001010"), -- i=1753
      ("10", "0111010111101110", "1110000000100100", "0110000000100100"), -- i=1754
      ("11", "0111010111101110", "1110000000100100", "1111010111101110"), -- i=1755
      ("00", "0001110011110011", "1110000110111000", "1111111010101011"), -- i=1756
      ("01", "0001110011110011", "1110000110111000", "0011101100111011"), -- i=1757
      ("10", "0001110011110011", "1110000110111000", "0000000010110000"), -- i=1758
      ("11", "0001110011110011", "1110000110111000", "1111110111111011"), -- i=1759
      ("00", "1101110001100011", "1001010001100001", "0111000011000100"), -- i=1760
      ("01", "1101110001100011", "1001010001100001", "0100100000000010"), -- i=1761
      ("10", "1101110001100011", "1001010001100001", "1001010001100001"), -- i=1762
      ("11", "1101110001100011", "1001010001100001", "1101110001100011"), -- i=1763
      ("00", "1000001110001110", "1010100011110101", "0010110010000011"), -- i=1764
      ("01", "1000001110001110", "1010100011110101", "1101101010011001"), -- i=1765
      ("10", "1000001110001110", "1010100011110101", "1000000010000100"), -- i=1766
      ("11", "1000001110001110", "1010100011110101", "1010101111111111"), -- i=1767
      ("00", "1010010101000111", "1110010101001011", "1000101010010010"), -- i=1768
      ("01", "1010010101000111", "1110010101001011", "1011111111111100"), -- i=1769
      ("10", "1010010101000111", "1110010101001011", "1010010101000011"), -- i=1770
      ("11", "1010010101000111", "1110010101001011", "1110010101001111"), -- i=1771
      ("00", "1100011011100100", "1100001110001011", "1000101001101111"), -- i=1772
      ("01", "1100011011100100", "1100001110001011", "0000001101011001"), -- i=1773
      ("10", "1100011011100100", "1100001110001011", "1100001010000000"), -- i=1774
      ("11", "1100011011100100", "1100001110001011", "1100011111101111"), -- i=1775
      ("00", "1101110111011100", "1100110010101101", "1010101010001001"), -- i=1776
      ("01", "1101110111011100", "1100110010101101", "0001000100101111"), -- i=1777
      ("10", "1101110111011100", "1100110010101101", "1100110010001100"), -- i=1778
      ("11", "1101110111011100", "1100110010101101", "1101110111111101"), -- i=1779
      ("00", "0001010111110101", "1000010111011000", "1001101111001101"), -- i=1780
      ("01", "0001010111110101", "1000010111011000", "1001000000011101"), -- i=1781
      ("10", "0001010111110101", "1000010111011000", "0000010111010000"), -- i=1782
      ("11", "0001010111110101", "1000010111011000", "1001010111111101"), -- i=1783
      ("00", "1111110011110101", "0000000010011111", "1111110110010100"), -- i=1784
      ("01", "1111110011110101", "0000000010011111", "1111110001010110"), -- i=1785
      ("10", "1111110011110101", "0000000010011111", "0000000010010101"), -- i=1786
      ("11", "1111110011110101", "0000000010011111", "1111110011111111"), -- i=1787
      ("00", "0110011111101101", "0101101001011010", "1100001001000111"), -- i=1788
      ("01", "0110011111101101", "0101101001011010", "0000110110010011"), -- i=1789
      ("10", "0110011111101101", "0101101001011010", "0100001001001000"), -- i=1790
      ("11", "0110011111101101", "0101101001011010", "0111111111111111"), -- i=1791
      ("00", "0101111011001011", "0100011011101110", "1010010110111001"), -- i=1792
      ("01", "0101111011001011", "0100011011101110", "0001011111011101"), -- i=1793
      ("10", "0101111011001011", "0100011011101110", "0100011011001010"), -- i=1794
      ("11", "0101111011001011", "0100011011101110", "0101111011101111"), -- i=1795
      ("00", "0101010111011011", "0110100111000010", "1011111110011101"), -- i=1796
      ("01", "0101010111011011", "0110100111000010", "1110110000011001"), -- i=1797
      ("10", "0101010111011011", "0110100111000010", "0100000111000010"), -- i=1798
      ("11", "0101010111011011", "0110100111000010", "0111110111011011"), -- i=1799
      ("00", "0000111111000111", "1111010000111010", "0000010000000001"), -- i=1800
      ("01", "0000111111000111", "1111010000111010", "0001101110001101"), -- i=1801
      ("10", "0000111111000111", "1111010000111010", "0000010000000010"), -- i=1802
      ("11", "0000111111000111", "1111010000111010", "1111111111111111"), -- i=1803
      ("00", "1101011010110010", "0010111010111001", "0000010101101011"), -- i=1804
      ("01", "1101011010110010", "0010111010111001", "1010011111111001"), -- i=1805
      ("10", "1101011010110010", "0010111010111001", "0000011010110000"), -- i=1806
      ("11", "1101011010110010", "0010111010111001", "1111111010111011"), -- i=1807
      ("00", "1100110100111011", "0001011101111111", "1110010010111010"), -- i=1808
      ("01", "1100110100111011", "0001011101111111", "1011010110111100"), -- i=1809
      ("10", "1100110100111011", "0001011101111111", "0000010100111011"), -- i=1810
      ("11", "1100110100111011", "0001011101111111", "1101111101111111"), -- i=1811
      ("00", "1111101000101111", "1011010001101100", "1010111010011011"), -- i=1812
      ("01", "1111101000101111", "1011010001101100", "0100010111000011"), -- i=1813
      ("10", "1111101000101111", "1011010001101100", "1011000000101100"), -- i=1814
      ("11", "1111101000101111", "1011010001101100", "1111111001101111"), -- i=1815
      ("00", "0100100001010100", "1001100110101110", "1110001000000010"), -- i=1816
      ("01", "0100100001010100", "1001100110101110", "1010111010100110"), -- i=1817
      ("10", "0100100001010100", "1001100110101110", "0000100000000100"), -- i=1818
      ("11", "0100100001010100", "1001100110101110", "1101100111111110"), -- i=1819
      ("00", "1111100010001011", "0011101001011010", "0011001011100101"), -- i=1820
      ("01", "1111100010001011", "0011101001011010", "1011111000110001"), -- i=1821
      ("10", "1111100010001011", "0011101001011010", "0011100000001010"), -- i=1822
      ("11", "1111100010001011", "0011101001011010", "1111101011011011"), -- i=1823
      ("00", "0100010010101010", "0000100001110010", "0100110100011100"), -- i=1824
      ("01", "0100010010101010", "0000100001110010", "0011110000111000"), -- i=1825
      ("10", "0100010010101010", "0000100001110010", "0000000000100010"), -- i=1826
      ("11", "0100010010101010", "0000100001110010", "0100110011111010"), -- i=1827
      ("00", "0000111000000011", "0001101100001001", "0010100100001100"), -- i=1828
      ("01", "0000111000000011", "0001101100001001", "1111001011111010"), -- i=1829
      ("10", "0000111000000011", "0001101100001001", "0000101000000001"), -- i=1830
      ("11", "0000111000000011", "0001101100001001", "0001111100001011"), -- i=1831
      ("00", "0010000100111101", "1101101001101101", "1111101110101010"), -- i=1832
      ("01", "0010000100111101", "1101101001101101", "0100011011010000"), -- i=1833
      ("10", "0010000100111101", "1101101001101101", "0000000000101101"), -- i=1834
      ("11", "0010000100111101", "1101101001101101", "1111101101111101"), -- i=1835
      ("00", "1010001010011001", "0001111010000100", "1100000100011101"), -- i=1836
      ("01", "1010001010011001", "0001111010000100", "1000010000010101"), -- i=1837
      ("10", "1010001010011001", "0001111010000100", "0000001010000000"), -- i=1838
      ("11", "1010001010011001", "0001111010000100", "1011111010011101"), -- i=1839
      ("00", "1011011111000001", "1011101001101100", "0111001000101101"), -- i=1840
      ("01", "1011011111000001", "1011101001101100", "1111110101010101"), -- i=1841
      ("10", "1011011111000001", "1011101001101100", "1011001001000000"), -- i=1842
      ("11", "1011011111000001", "1011101001101100", "1011111111101101"), -- i=1843
      ("00", "0010111110101011", "1101010011011101", "0000010010001000"), -- i=1844
      ("01", "0010111110101011", "1101010011011101", "0101101011001110"), -- i=1845
      ("10", "0010111110101011", "1101010011011101", "0000010010001001"), -- i=1846
      ("11", "0010111110101011", "1101010011011101", "1111111111111111"), -- i=1847
      ("00", "0100001110001111", "1100111001100010", "0001000111110001"), -- i=1848
      ("01", "0100001110001111", "1100111001100010", "0111010100101101"), -- i=1849
      ("10", "0100001110001111", "1100111001100010", "0100001000000010"), -- i=1850
      ("11", "0100001110001111", "1100111001100010", "1100111111101111"), -- i=1851
      ("00", "0010111000101111", "0011000000000101", "0101111000110100"), -- i=1852
      ("01", "0010111000101111", "0011000000000101", "1111111000101010"), -- i=1853
      ("10", "0010111000101111", "0011000000000101", "0010000000000101"), -- i=1854
      ("11", "0010111000101111", "0011000000000101", "0011111000101111"), -- i=1855
      ("00", "0010111010011001", "1111111000111100", "0010110011010101"), -- i=1856
      ("01", "0010111010011001", "1111111000111100", "0011000001011101"), -- i=1857
      ("10", "0010111010011001", "1111111000111100", "0010111000011000"), -- i=1858
      ("11", "0010111010011001", "1111111000111100", "1111111010111101"), -- i=1859
      ("00", "0001100110110110", "0101011111000011", "0111000101111001"), -- i=1860
      ("01", "0001100110110110", "0101011111000011", "1100000111110011"), -- i=1861
      ("10", "0001100110110110", "0101011111000011", "0001000110000010"), -- i=1862
      ("11", "0001100110110110", "0101011111000011", "0101111111110111"), -- i=1863
      ("00", "0011100000110100", "1111010111000000", "0010110111110100"), -- i=1864
      ("01", "0011100000110100", "1111010111000000", "0100001001110100"), -- i=1865
      ("10", "0011100000110100", "1111010111000000", "0011000000000000"), -- i=1866
      ("11", "0011100000110100", "1111010111000000", "1111110111110100"), -- i=1867
      ("00", "0011110110010010", "1001110110010011", "1101101100100101"), -- i=1868
      ("01", "0011110110010010", "1001110110010011", "1001111111111111"), -- i=1869
      ("10", "0011110110010010", "1001110110010011", "0001110110010010"), -- i=1870
      ("11", "0011110110010010", "1001110110010011", "1011110110010011"), -- i=1871
      ("00", "0110011010011010", "1111110000100100", "0110001010111110"), -- i=1872
      ("01", "0110011010011010", "1111110000100100", "0110101001110110"), -- i=1873
      ("10", "0110011010011010", "1111110000100100", "0110010000000000"), -- i=1874
      ("11", "0110011010011010", "1111110000100100", "1111111010111110"), -- i=1875
      ("00", "1001001010110001", "1000100110101111", "0001110001100000"), -- i=1876
      ("01", "1001001010110001", "1000100110101111", "0000100100000010"), -- i=1877
      ("10", "1001001010110001", "1000100110101111", "1000000010100001"), -- i=1878
      ("11", "1001001010110001", "1000100110101111", "1001101110111111"), -- i=1879
      ("00", "1001100101110111", "1100001100000100", "0101110001111011"), -- i=1880
      ("01", "1001100101110111", "1100001100000100", "1101011001110011"), -- i=1881
      ("10", "1001100101110111", "1100001100000100", "1000000100000100"), -- i=1882
      ("11", "1001100101110111", "1100001100000100", "1101101101110111"), -- i=1883
      ("00", "0110111000001110", "0011010110100101", "1010001110110011"), -- i=1884
      ("01", "0110111000001110", "0011010110100101", "0011100001101001"), -- i=1885
      ("10", "0110111000001110", "0011010110100101", "0010010000000100"), -- i=1886
      ("11", "0110111000001110", "0011010110100101", "0111111110101111"), -- i=1887
      ("00", "0110000011100110", "1111110111010110", "0101111010111100"), -- i=1888
      ("01", "0110000011100110", "1111110111010110", "0110001100010000"), -- i=1889
      ("10", "0110000011100110", "1111110111010110", "0110000011000110"), -- i=1890
      ("11", "0110000011100110", "1111110111010110", "1111110111110110"), -- i=1891
      ("00", "0010000011001010", "1000110000011100", "1010110011100110"), -- i=1892
      ("01", "0010000011001010", "1000110000011100", "1001010010101110"), -- i=1893
      ("10", "0010000011001010", "1000110000011100", "0000000000001000"), -- i=1894
      ("11", "0010000011001010", "1000110000011100", "1010110011011110"), -- i=1895
      ("00", "1111000110100010", "1110101000101001", "1101101111001011"), -- i=1896
      ("01", "1111000110100010", "1110101000101001", "0000011101111001"), -- i=1897
      ("10", "1111000110100010", "1110101000101001", "1110000000100000"), -- i=1898
      ("11", "1111000110100010", "1110101000101001", "1111101110101011"), -- i=1899
      ("00", "1111010001011000", "1001000010111111", "1000010100010111"), -- i=1900
      ("01", "1111010001011000", "1001000010111111", "0110001110011001"), -- i=1901
      ("10", "1111010001011000", "1001000010111111", "1001000000011000"), -- i=1902
      ("11", "1111010001011000", "1001000010111111", "1111010011111111"), -- i=1903
      ("00", "1010110001100011", "1111000000100000", "1001110010000011"), -- i=1904
      ("01", "1010110001100011", "1111000000100000", "1011110001000011"), -- i=1905
      ("10", "1010110001100011", "1111000000100000", "1010000000100000"), -- i=1906
      ("11", "1010110001100011", "1111000000100000", "1111110001100011"), -- i=1907
      ("00", "0001111000111100", "1000011001110000", "1010010010101100"), -- i=1908
      ("01", "0001111000111100", "1000011001110000", "1001011111001100"), -- i=1909
      ("10", "0001111000111100", "1000011001110000", "0000011000110000"), -- i=1910
      ("11", "0001111000111100", "1000011001110000", "1001111001111100"), -- i=1911
      ("00", "1011001110100110", "0010101000010110", "1101110110111100"), -- i=1912
      ("01", "1011001110100110", "0010101000010110", "1000100110010000"), -- i=1913
      ("10", "1011001110100110", "0010101000010110", "0010001000000110"), -- i=1914
      ("11", "1011001110100110", "0010101000010110", "1011101110110110"), -- i=1915
      ("00", "0110000001001111", "1010010100101110", "0000010101111101"), -- i=1916
      ("01", "0110000001001111", "1010010100101110", "1011101100100001"), -- i=1917
      ("10", "0110000001001111", "1010010100101110", "0010000000001110"), -- i=1918
      ("11", "0110000001001111", "1010010100101110", "1110010101101111"), -- i=1919
      ("00", "0111100001001101", "1111000101010101", "0110100110100010"), -- i=1920
      ("01", "0111100001001101", "1111000101010101", "1000011011111000"), -- i=1921
      ("10", "0111100001001101", "1111000101010101", "0111000001000101"), -- i=1922
      ("11", "0111100001001101", "1111000101010101", "1111100101011101"), -- i=1923
      ("00", "0000101110010110", "0001010001011010", "0001111111110000"), -- i=1924
      ("01", "0000101110010110", "0001010001011010", "1111011100111100"), -- i=1925
      ("10", "0000101110010110", "0001010001011010", "0000000000010010"), -- i=1926
      ("11", "0000101110010110", "0001010001011010", "0001111111011110"), -- i=1927
      ("00", "1111101011100010", "1000010100111101", "1000000000011111"), -- i=1928
      ("01", "1111101011100010", "1000010100111101", "0111010110100101"), -- i=1929
      ("10", "1111101011100010", "1000010100111101", "1000000000100000"), -- i=1930
      ("11", "1111101011100010", "1000010100111101", "1111111111111111"), -- i=1931
      ("00", "0000010100000101", "0000100101000000", "0000111001000101"), -- i=1932
      ("01", "0000010100000101", "0000100101000000", "1111101111000101"), -- i=1933
      ("10", "0000010100000101", "0000100101000000", "0000000100000000"), -- i=1934
      ("11", "0000010100000101", "0000100101000000", "0000110101000101"), -- i=1935
      ("00", "1011110001100110", "1000000101100011", "0011110111001001"), -- i=1936
      ("01", "1011110001100110", "1000000101100011", "0011101100000011"), -- i=1937
      ("10", "1011110001100110", "1000000101100011", "1000000001100010"), -- i=1938
      ("11", "1011110001100110", "1000000101100011", "1011110101100111"), -- i=1939
      ("00", "0011110011010011", "0011110100011011", "0111100111101110"), -- i=1940
      ("01", "0011110011010011", "0011110100011011", "1111111110111000"), -- i=1941
      ("10", "0011110011010011", "0011110100011011", "0011110000010011"), -- i=1942
      ("11", "0011110011010011", "0011110100011011", "0011110111011011"), -- i=1943
      ("00", "1111111011110110", "0001111001101000", "0001110101011110"), -- i=1944
      ("01", "1111111011110110", "0001111001101000", "1110000010001110"), -- i=1945
      ("10", "1111111011110110", "0001111001101000", "0001111001100000"), -- i=1946
      ("11", "1111111011110110", "0001111001101000", "1111111011111110"), -- i=1947
      ("00", "1100001000100110", "0110100011101000", "0010101100001110"), -- i=1948
      ("01", "1100001000100110", "0110100011101000", "0101100100111110"), -- i=1949
      ("10", "1100001000100110", "0110100011101000", "0100000000100000"), -- i=1950
      ("11", "1100001000100110", "0110100011101000", "1110101011101110"), -- i=1951
      ("00", "0000001110110011", "0010100010011111", "0010110001010010"), -- i=1952
      ("01", "0000001110110011", "0010100010011111", "1101101100010100"), -- i=1953
      ("10", "0000001110110011", "0010100010011111", "0000000010010011"), -- i=1954
      ("11", "0000001110110011", "0010100010011111", "0010101110111111"), -- i=1955
      ("00", "0011111001000111", "0001100011001010", "0101011100010001"), -- i=1956
      ("01", "0011111001000111", "0001100011001010", "0010010101111101"), -- i=1957
      ("10", "0011111001000111", "0001100011001010", "0001100001000010"), -- i=1958
      ("11", "0011111001000111", "0001100011001010", "0011111011001111"), -- i=1959
      ("00", "0110100010101110", "0010111011000011", "1001011101110001"), -- i=1960
      ("01", "0110100010101110", "0010111011000011", "0011100111101011"), -- i=1961
      ("10", "0110100010101110", "0010111011000011", "0010100010000010"), -- i=1962
      ("11", "0110100010101110", "0010111011000011", "0110111011101111"), -- i=1963
      ("00", "0010101110101011", "1111001111011000", "0001111110000011"), -- i=1964
      ("01", "0010101110101011", "1111001111011000", "0011011111010011"), -- i=1965
      ("10", "0010101110101011", "1111001111011000", "0010001110001000"), -- i=1966
      ("11", "0010101110101011", "1111001111011000", "1111101111111011"), -- i=1967
      ("00", "1010011011010001", "1010101001001000", "0101000100011001"), -- i=1968
      ("01", "1010011011010001", "1010101001001000", "1111110010001001"), -- i=1969
      ("10", "1010011011010001", "1010101001001000", "1010001001000000"), -- i=1970
      ("11", "1010011011010001", "1010101001001000", "1010111011011001"), -- i=1971
      ("00", "1000111001100011", "1000100010001000", "0001011011101011"), -- i=1972
      ("01", "1000111001100011", "1000100010001000", "0000010111011011"), -- i=1973
      ("10", "1000111001100011", "1000100010001000", "1000100000000000"), -- i=1974
      ("11", "1000111001100011", "1000100010001000", "1000111011101011"), -- i=1975
      ("00", "1111010011111111", "1100101000010110", "1011111100010101"), -- i=1976
      ("01", "1111010011111111", "1100101000010110", "0010101011101001"), -- i=1977
      ("10", "1111010011111111", "1100101000010110", "1100000000010110"), -- i=1978
      ("11", "1111010011111111", "1100101000010110", "1111111011111111"), -- i=1979
      ("00", "0100110011101001", "1100100100010110", "0001010111111111"), -- i=1980
      ("01", "0100110011101001", "1100100100010110", "1000001111010011"), -- i=1981
      ("10", "0100110011101001", "1100100100010110", "0100100000000000"), -- i=1982
      ("11", "0100110011101001", "1100100100010110", "1100110111111111"), -- i=1983
      ("00", "1000001011011110", "0001011110110111", "1001101010010101"), -- i=1984
      ("01", "1000001011011110", "0001011110110111", "0110101100100111"), -- i=1985
      ("10", "1000001011011110", "0001011110110111", "0000001010010110"), -- i=1986
      ("11", "1000001011011110", "0001011110110111", "1001011111111111"), -- i=1987
      ("00", "1000100101000011", "1010011010101001", "0010111111101100"), -- i=1988
      ("01", "1000100101000011", "1010011010101001", "1110001010011010"), -- i=1989
      ("10", "1000100101000011", "1010011010101001", "1000000000000001"), -- i=1990
      ("11", "1000100101000011", "1010011010101001", "1010111111101011"), -- i=1991
      ("00", "0001001100011000", "0110011000110101", "0111100101001101"), -- i=1992
      ("01", "0001001100011000", "0110011000110101", "1010110011100011"), -- i=1993
      ("10", "0001001100011000", "0110011000110101", "0000001000010000"), -- i=1994
      ("11", "0001001100011000", "0110011000110101", "0111011100111101"), -- i=1995
      ("00", "1000001111101101", "1010010011111010", "0010100011100111"), -- i=1996
      ("01", "1000001111101101", "1010010011111010", "1101111011110011"), -- i=1997
      ("10", "1000001111101101", "1010010011111010", "1000000011101000"), -- i=1998
      ("11", "1000001111101101", "1010010011111010", "1010011111111111"), -- i=1999
      ("00", "0111100111110011", "0101100101001011", "1101001100111110"), -- i=2000
      ("01", "0111100111110011", "0101100101001011", "0010000010101000"), -- i=2001
      ("10", "0111100111110011", "0101100101001011", "0101100101000011"), -- i=2002
      ("11", "0111100111110011", "0101100101001011", "0111100111111011"), -- i=2003
      ("00", "1010001100011100", "1101001111010010", "0111011011101110"), -- i=2004
      ("01", "1010001100011100", "1101001111010010", "1100111101001010"), -- i=2005
      ("10", "1010001100011100", "1101001111010010", "1000001100010000"), -- i=2006
      ("11", "1010001100011100", "1101001111010010", "1111001111011110"), -- i=2007
      ("00", "0110101010001100", "0101101010011101", "1100010100101001"), -- i=2008
      ("01", "0110101010001100", "0101101010011101", "0000111111101111"), -- i=2009
      ("10", "0110101010001100", "0101101010011101", "0100101010001100"), -- i=2010
      ("11", "0110101010001100", "0101101010011101", "0111101010011101"), -- i=2011
      ("00", "0011001000110000", "0101011010100110", "1000100011010110"), -- i=2012
      ("01", "0011001000110000", "0101011010100110", "1101101110001010"), -- i=2013
      ("10", "0011001000110000", "0101011010100110", "0001001000100000"), -- i=2014
      ("11", "0011001000110000", "0101011010100110", "0111011010110110"), -- i=2015
      ("00", "0100101000110010", "0000001000000101", "0100110000110111"), -- i=2016
      ("01", "0100101000110010", "0000001000000101", "0100100000101101"), -- i=2017
      ("10", "0100101000110010", "0000001000000101", "0000001000000000"), -- i=2018
      ("11", "0100101000110010", "0000001000000101", "0100101000110111"), -- i=2019
      ("00", "0100111001111000", "1000011000001100", "1101010010000100"), -- i=2020
      ("01", "0100111001111000", "1000011000001100", "1100100001101100"), -- i=2021
      ("10", "0100111001111000", "1000011000001100", "0000011000001000"), -- i=2022
      ("11", "0100111001111000", "1000011000001100", "1100111001111100"), -- i=2023
      ("00", "0111011010000110", "1100110101010000", "0100001111010110"), -- i=2024
      ("01", "0111011010000110", "1100110101010000", "1010100100110110"), -- i=2025
      ("10", "0111011010000110", "1100110101010000", "0100010000000000"), -- i=2026
      ("11", "0111011010000110", "1100110101010000", "1111111111010110"), -- i=2027
      ("00", "0011111110011100", "1100000111110011", "0000000110001111"), -- i=2028
      ("01", "0011111110011100", "1100000111110011", "0111110110101001"), -- i=2029
      ("10", "0011111110011100", "1100000111110011", "0000000110010000"), -- i=2030
      ("11", "0011111110011100", "1100000111110011", "1111111111111111"), -- i=2031
      ("00", "1000100001110001", "1000001011010110", "0000101101000111"), -- i=2032
      ("01", "1000100001110001", "1000001011010110", "0000010110011011"), -- i=2033
      ("10", "1000100001110001", "1000001011010110", "1000000001010000"), -- i=2034
      ("11", "1000100001110001", "1000001011010110", "1000101011110111"), -- i=2035
      ("00", "0010101101000110", "0011111011000101", "0110101000001011"), -- i=2036
      ("01", "0010101101000110", "0011111011000101", "1110110010000001"), -- i=2037
      ("10", "0010101101000110", "0011111011000101", "0010101001000100"), -- i=2038
      ("11", "0010101101000110", "0011111011000101", "0011111111000111"), -- i=2039
      ("00", "1010001100011011", "1100000111011100", "0110010011110111"), -- i=2040
      ("01", "1010001100011011", "1100000111011100", "1110000100111111"), -- i=2041
      ("10", "1010001100011011", "1100000111011100", "1000000100011000"), -- i=2042
      ("11", "1010001100011011", "1100000111011100", "1110001111011111"), -- i=2043
      ("00", "1010110011101010", "0111001011010010", "0001111110111100"), -- i=2044
      ("01", "1010110011101010", "0111001011010010", "0011101000011000"), -- i=2045
      ("10", "1010110011101010", "0111001011010010", "0010000011000010"), -- i=2046
      ("11", "1010110011101010", "0111001011010010", "1111111011111010"), -- i=2047
      ("00", "1100101101101000", "0001001010100101", "1101111000001101"), -- i=2048
      ("01", "1100101101101000", "0001001010100101", "1011100011000011"), -- i=2049
      ("10", "1100101101101000", "0001001010100101", "0000001000100000"), -- i=2050
      ("11", "1100101101101000", "0001001010100101", "1101101111101101"), -- i=2051
      ("00", "0101101111000000", "0100110011001101", "1010100010001101"), -- i=2052
      ("01", "0101101111000000", "0100110011001101", "0000111011110011"), -- i=2053
      ("10", "0101101111000000", "0100110011001101", "0100100011000000"), -- i=2054
      ("11", "0101101111000000", "0100110011001101", "0101111111001101"), -- i=2055
      ("00", "1001100110101010", "0011111110011011", "1101100101000101"), -- i=2056
      ("01", "1001100110101010", "0011111110011011", "0101101000001111"), -- i=2057
      ("10", "1001100110101010", "0011111110011011", "0001100110001010"), -- i=2058
      ("11", "1001100110101010", "0011111110011011", "1011111110111011"), -- i=2059
      ("00", "1011001001001110", "0000011100011011", "1011100101101001"), -- i=2060
      ("01", "1011001001001110", "0000011100011011", "1010101100110011"), -- i=2061
      ("10", "1011001001001110", "0000011100011011", "0000001000001010"), -- i=2062
      ("11", "1011001001001110", "0000011100011011", "1011011101011111"), -- i=2063
      ("00", "0101010010000110", "1110000000000110", "0011010010001100"), -- i=2064
      ("01", "0101010010000110", "1110000000000110", "0111010010000000"), -- i=2065
      ("10", "0101010010000110", "1110000000000110", "0100000000000110"), -- i=2066
      ("11", "0101010010000110", "1110000000000110", "1111010010000110"), -- i=2067
      ("00", "0001110000100000", "0011111101000011", "0101101101100011"), -- i=2068
      ("01", "0001110000100000", "0011111101000011", "1101110011011101"), -- i=2069
      ("10", "0001110000100000", "0011111101000011", "0001110000000000"), -- i=2070
      ("11", "0001110000100000", "0011111101000011", "0011111101100011"), -- i=2071
      ("00", "1010100101010010", "1100010000100100", "0110110101110110"), -- i=2072
      ("01", "1010100101010010", "1100010000100100", "1110010100101110"), -- i=2073
      ("10", "1010100101010010", "1100010000100100", "1000000000000000"), -- i=2074
      ("11", "1010100101010010", "1100010000100100", "1110110101110110"), -- i=2075
      ("00", "0010011101111011", "1111001111010101", "0001101101010000"), -- i=2076
      ("01", "0010011101111011", "1111001111010101", "0011001110100110"), -- i=2077
      ("10", "0010011101111011", "1111001111010101", "0010001101010001"), -- i=2078
      ("11", "0010011101111011", "1111001111010101", "1111011111111111"), -- i=2079
      ("00", "1100001101001010", "0110000110101010", "0010010011110100"), -- i=2080
      ("01", "1100001101001010", "0110000110101010", "0110000110100000"), -- i=2081
      ("10", "1100001101001010", "0110000110101010", "0100000100001010"), -- i=2082
      ("11", "1100001101001010", "0110000110101010", "1110001111101010"), -- i=2083
      ("00", "1111101000110011", "0010111001110100", "0010100010100111"), -- i=2084
      ("01", "1111101000110011", "0010111001110100", "1100101110111111"), -- i=2085
      ("10", "1111101000110011", "0010111001110100", "0010101000110000"), -- i=2086
      ("11", "1111101000110011", "0010111001110100", "1111111001110111"), -- i=2087
      ("00", "0111100001111100", "0111011011110011", "1110111101101111"), -- i=2088
      ("01", "0111100001111100", "0111011011110011", "0000000110001001"), -- i=2089
      ("10", "0111100001111100", "0111011011110011", "0111000001110000"), -- i=2090
      ("11", "0111100001111100", "0111011011110011", "0111111011111111"), -- i=2091
      ("00", "0011000111111001", "0110101011110101", "1001110011101110"), -- i=2092
      ("01", "0011000111111001", "0110101011110101", "1100011100000100"), -- i=2093
      ("10", "0011000111111001", "0110101011110101", "0010000011110001"), -- i=2094
      ("11", "0011000111111001", "0110101011110101", "0111101111111101"), -- i=2095
      ("00", "1010000000111011", "1101101001111000", "0111101010110011"), -- i=2096
      ("01", "1010000000111011", "1101101001111000", "1100010111000011"), -- i=2097
      ("10", "1010000000111011", "1101101001111000", "1000000000111000"), -- i=2098
      ("11", "1010000000111011", "1101101001111000", "1111101001111011"), -- i=2099
      ("00", "0100100110110101", "0011111110110011", "1000100101101000"), -- i=2100
      ("01", "0100100110110101", "0011111110110011", "0000101000000010"), -- i=2101
      ("10", "0100100110110101", "0011111110110011", "0000100110110001"), -- i=2102
      ("11", "0100100110110101", "0011111110110011", "0111111110110111"), -- i=2103
      ("00", "0110110001111010", "1101001101000001", "0011111110111011"), -- i=2104
      ("01", "0110110001111010", "1101001101000001", "1001100100111001"), -- i=2105
      ("10", "0110110001111010", "1101001101000001", "0100000001000000"), -- i=2106
      ("11", "0110110001111010", "1101001101000001", "1111111101111011"), -- i=2107
      ("00", "0111011011010001", "0110011010001010", "1101110101011011"), -- i=2108
      ("01", "0111011011010001", "0110011010001010", "0001000001000111"), -- i=2109
      ("10", "0111011011010001", "0110011010001010", "0110011010000000"), -- i=2110
      ("11", "0111011011010001", "0110011010001010", "0111011011011011"), -- i=2111
      ("00", "1100110001101101", "0110011001101100", "0011001011011001"), -- i=2112
      ("01", "1100110001101101", "0110011001101100", "0110011000000001"), -- i=2113
      ("10", "1100110001101101", "0110011001101100", "0100010001101100"), -- i=2114
      ("11", "1100110001101101", "0110011001101100", "1110111001101101"), -- i=2115
      ("00", "1011001010000111", "0000100100100000", "1011101110100111"), -- i=2116
      ("01", "1011001010000111", "0000100100100000", "1010100101100111"), -- i=2117
      ("10", "1011001010000111", "0000100100100000", "0000000000000000"), -- i=2118
      ("11", "1011001010000111", "0000100100100000", "1011101110100111"), -- i=2119
      ("00", "0111010000110111", "1011110100010011", "0011000101001010"), -- i=2120
      ("01", "0111010000110111", "1011110100010011", "1011011100100100"), -- i=2121
      ("10", "0111010000110111", "1011110100010011", "0011010000010011"), -- i=2122
      ("11", "0111010000110111", "1011110100010011", "1111110100110111"), -- i=2123
      ("00", "0100110010001100", "0001111001100010", "0110101011101110"), -- i=2124
      ("01", "0100110010001100", "0001111001100010", "0010111000101010"), -- i=2125
      ("10", "0100110010001100", "0001111001100010", "0000110000000000"), -- i=2126
      ("11", "0100110010001100", "0001111001100010", "0101111011101110"), -- i=2127
      ("00", "0010001010011110", "0010010100010011", "0100011110110001"), -- i=2128
      ("01", "0010001010011110", "0010010100010011", "1111110110001011"), -- i=2129
      ("10", "0010001010011110", "0010010100010011", "0010000000010010"), -- i=2130
      ("11", "0010001010011110", "0010010100010011", "0010011110011111"), -- i=2131
      ("00", "1111010110111010", "1011101001100111", "1011000000100001"), -- i=2132
      ("01", "1111010110111010", "1011101001100111", "0011101101010011"), -- i=2133
      ("10", "1111010110111010", "1011101001100111", "1011000000100010"), -- i=2134
      ("11", "1111010110111010", "1011101001100111", "1111111111111111"), -- i=2135
      ("00", "0010001011111100", "0011011001111111", "0101100101111011"), -- i=2136
      ("01", "0010001011111100", "0011011001111111", "1110110001111101"), -- i=2137
      ("10", "0010001011111100", "0011011001111111", "0010001001111100"), -- i=2138
      ("11", "0010001011111100", "0011011001111111", "0011011011111111"), -- i=2139
      ("00", "1010101010000101", "0110110100011111", "0001011110100100"), -- i=2140
      ("01", "1010101010000101", "0110110100011111", "0011110101100110"), -- i=2141
      ("10", "1010101010000101", "0110110100011111", "0010100000000101"), -- i=2142
      ("11", "1010101010000101", "0110110100011111", "1110111110011111"), -- i=2143
      ("00", "1101011011101000", "0101011011010011", "0010110110111011"), -- i=2144
      ("01", "1101011011101000", "0101011011010011", "1000000000010101"), -- i=2145
      ("10", "1101011011101000", "0101011011010011", "0101011011000000"), -- i=2146
      ("11", "1101011011101000", "0101011011010011", "1101011011111011"), -- i=2147
      ("00", "0100011001100111", "0010111101110001", "0111010111011000"), -- i=2148
      ("01", "0100011001100111", "0010111101110001", "0001011011110110"), -- i=2149
      ("10", "0100011001100111", "0010111101110001", "0000011001100001"), -- i=2150
      ("11", "0100011001100111", "0010111101110001", "0110111101110111"), -- i=2151
      ("00", "0100100001001111", "0010101000100000", "0111001001101111"), -- i=2152
      ("01", "0100100001001111", "0010101000100000", "0001111000101111"), -- i=2153
      ("10", "0100100001001111", "0010101000100000", "0000100000000000"), -- i=2154
      ("11", "0100100001001111", "0010101000100000", "0110101001101111"), -- i=2155
      ("00", "1101001010001110", "1110100111000101", "1011110001010011"), -- i=2156
      ("01", "1101001010001110", "1110100111000101", "1110100011001001"), -- i=2157
      ("10", "1101001010001110", "1110100111000101", "1100000010000100"), -- i=2158
      ("11", "1101001010001110", "1110100111000101", "1111101111001111"), -- i=2159
      ("00", "0110001000000000", "1000000111010001", "1110001111010001"), -- i=2160
      ("01", "0110001000000000", "1000000111010001", "1110000000101111"), -- i=2161
      ("10", "0110001000000000", "1000000111010001", "0000000000000000"), -- i=2162
      ("11", "0110001000000000", "1000000111010001", "1110001111010001"), -- i=2163
      ("00", "1101001101100111", "0101001000001001", "0010010101110000"), -- i=2164
      ("01", "1101001101100111", "0101001000001001", "1000000101011110"), -- i=2165
      ("10", "1101001101100111", "0101001000001001", "0101001000000001"), -- i=2166
      ("11", "1101001101100111", "0101001000001001", "1101001101101111"), -- i=2167
      ("00", "0111000111011000", "1111111110111101", "0111000110010101"), -- i=2168
      ("01", "0111000111011000", "1111111110111101", "0111001000011011"), -- i=2169
      ("10", "0111000111011000", "1111111110111101", "0111000110011000"), -- i=2170
      ("11", "0111000111011000", "1111111110111101", "1111111111111101"), -- i=2171
      ("00", "1111000111101110", "1011101010111000", "1010110010100110"), -- i=2172
      ("01", "1111000111101110", "1011101010111000", "0011011100110110"), -- i=2173
      ("10", "1111000111101110", "1011101010111000", "1011000010101000"), -- i=2174
      ("11", "1111000111101110", "1011101010111000", "1111101111111110"), -- i=2175
      ("00", "0000010100010010", "1111001110011110", "1111100010110000"), -- i=2176
      ("01", "0000010100010010", "1111001110011110", "0001000101110100"), -- i=2177
      ("10", "0000010100010010", "1111001110011110", "0000000100010010"), -- i=2178
      ("11", "0000010100010010", "1111001110011110", "1111011110011110"), -- i=2179
      ("00", "0101111011001110", "0110111101110101", "1100111001000011"), -- i=2180
      ("01", "0101111011001110", "0110111101110101", "1110111101011001"), -- i=2181
      ("10", "0101111011001110", "0110111101110101", "0100111001000100"), -- i=2182
      ("11", "0101111011001110", "0110111101110101", "0111111111111111"), -- i=2183
      ("00", "0000010001101101", "1111000000101111", "1111010010011100"), -- i=2184
      ("01", "0000010001101101", "1111000000101111", "0001010000111110"), -- i=2185
      ("10", "0000010001101101", "1111000000101111", "0000000000101101"), -- i=2186
      ("11", "0000010001101101", "1111000000101111", "1111010001101111"), -- i=2187
      ("00", "0011011010101111", "0110011100110000", "1001110111011111"), -- i=2188
      ("01", "0011011010101111", "0110011100110000", "1100111101111111"), -- i=2189
      ("10", "0011011010101111", "0110011100110000", "0010011000100000"), -- i=2190
      ("11", "0011011010101111", "0110011100110000", "0111011110111111"), -- i=2191
      ("00", "0011001100101100", "0011010010001001", "0110011110110101"), -- i=2192
      ("01", "0011001100101100", "0011010010001001", "1111111010100011"), -- i=2193
      ("10", "0011001100101100", "0011010010001001", "0011000000001000"), -- i=2194
      ("11", "0011001100101100", "0011010010001001", "0011011110101101"), -- i=2195
      ("00", "0000000001001111", "0110011100000011", "0110011101010010"), -- i=2196
      ("01", "0000000001001111", "0110011100000011", "1001100101001100"), -- i=2197
      ("10", "0000000001001111", "0110011100000011", "0000000000000011"), -- i=2198
      ("11", "0000000001001111", "0110011100000011", "0110011101001111"), -- i=2199
      ("00", "1101100100011111", "0100110101101110", "0010011010001101"), -- i=2200
      ("01", "1101100100011111", "0100110101101110", "1000101110110001"), -- i=2201
      ("10", "1101100100011111", "0100110101101110", "0100100100001110"), -- i=2202
      ("11", "1101100100011111", "0100110101101110", "1101110101111111"), -- i=2203
      ("00", "0001011000111111", "0010110000100000", "0100001001011111"), -- i=2204
      ("01", "0001011000111111", "0010110000100000", "1110101000011111"), -- i=2205
      ("10", "0001011000111111", "0010110000100000", "0000010000100000"), -- i=2206
      ("11", "0001011000111111", "0010110000100000", "0011111000111111"), -- i=2207
      ("00", "0110110100111011", "0100000110101111", "1010111011101010"), -- i=2208
      ("01", "0110110100111011", "0100000110101111", "0010101110001100"), -- i=2209
      ("10", "0110110100111011", "0100000110101111", "0100000100101011"), -- i=2210
      ("11", "0110110100111011", "0100000110101111", "0110110110111111"), -- i=2211
      ("00", "0110111101011111", "1101011010001101", "0100010111101100"), -- i=2212
      ("01", "0110111101011111", "1101011010001101", "1001100011010010"), -- i=2213
      ("10", "0110111101011111", "1101011010001101", "0100011000001101"), -- i=2214
      ("11", "0110111101011111", "1101011010001101", "1111111111011111"), -- i=2215
      ("00", "1000101101101010", "0011001111010111", "1011111101000001"), -- i=2216
      ("01", "1000101101101010", "0011001111010111", "0101011110010011"), -- i=2217
      ("10", "1000101101101010", "0011001111010111", "0000001101000010"), -- i=2218
      ("11", "1000101101101010", "0011001111010111", "1011101111111111"), -- i=2219
      ("00", "1100001001101010", "1001100110001111", "0101101111111001"), -- i=2220
      ("01", "1100001001101010", "1001100110001111", "0010100011011011"), -- i=2221
      ("10", "1100001001101010", "1001100110001111", "1000000000001010"), -- i=2222
      ("11", "1100001001101010", "1001100110001111", "1101101111101111"), -- i=2223
      ("00", "0101110110100011", "1010001010111010", "0000000001011101"), -- i=2224
      ("01", "0101110110100011", "1010001010111010", "1011101011101001"), -- i=2225
      ("10", "0101110110100011", "1010001010111010", "0000000010100010"), -- i=2226
      ("11", "0101110110100011", "1010001010111010", "1111111110111011"), -- i=2227
      ("00", "0111001000111101", "1010100111101010", "0001110000100111"), -- i=2228
      ("01", "0111001000111101", "1010100111101010", "1100100001010011"), -- i=2229
      ("10", "0111001000111101", "1010100111101010", "0010000000101000"), -- i=2230
      ("11", "0111001000111101", "1010100111101010", "1111101111111111"), -- i=2231
      ("00", "1110010101101111", "0101100110101001", "0011111100011000"), -- i=2232
      ("01", "1110010101101111", "0101100110101001", "1000101111000110"), -- i=2233
      ("10", "1110010101101111", "0101100110101001", "0100000100101001"), -- i=2234
      ("11", "1110010101101111", "0101100110101001", "1111110111101111"), -- i=2235
      ("00", "0000100110100010", "0111110101101011", "1000011100001101"), -- i=2236
      ("01", "0000100110100010", "0111110101101011", "1000110000110111"), -- i=2237
      ("10", "0000100110100010", "0111110101101011", "0000100100100010"), -- i=2238
      ("11", "0000100110100010", "0111110101101011", "0111110111101011"), -- i=2239
      ("00", "0100000001100100", "1011000001010101", "1111000010111001"), -- i=2240
      ("01", "0100000001100100", "1011000001010101", "1001000000001111"), -- i=2241
      ("10", "0100000001100100", "1011000001010101", "0000000001000100"), -- i=2242
      ("11", "0100000001100100", "1011000001010101", "1111000001110101"), -- i=2243
      ("00", "0100111011000010", "1011001001011011", "0000000100011101"), -- i=2244
      ("01", "0100111011000010", "1011001001011011", "1001110001100111"), -- i=2245
      ("10", "0100111011000010", "1011001001011011", "0000001001000010"), -- i=2246
      ("11", "0100111011000010", "1011001001011011", "1111111011011011"), -- i=2247
      ("00", "0001011101000111", "1111000110110001", "0000100011111000"), -- i=2248
      ("01", "0001011101000111", "1111000110110001", "0010010110010110"), -- i=2249
      ("10", "0001011101000111", "1111000110110001", "0001000100000001"), -- i=2250
      ("11", "0001011101000111", "1111000110110001", "1111011111110111"), -- i=2251
      ("00", "0001111110011101", "0110000011001100", "1000000001101001"), -- i=2252
      ("01", "0001111110011101", "0110000011001100", "1011111011010001"), -- i=2253
      ("10", "0001111110011101", "0110000011001100", "0000000010001100"), -- i=2254
      ("11", "0001111110011101", "0110000011001100", "0111111111011101"), -- i=2255
      ("00", "1110010011010110", "1010000001010101", "1000010100101011"), -- i=2256
      ("01", "1110010011010110", "1010000001010101", "0100010010000001"), -- i=2257
      ("10", "1110010011010110", "1010000001010101", "1010000001010100"), -- i=2258
      ("11", "1110010011010110", "1010000001010101", "1110010011010111"), -- i=2259
      ("00", "0101101000001101", "0010101011100111", "1000010011110100"), -- i=2260
      ("01", "0101101000001101", "0010101011100111", "0010111100100110"), -- i=2261
      ("10", "0101101000001101", "0010101011100111", "0000101000000101"), -- i=2262
      ("11", "0101101000001101", "0010101011100111", "0111101011101111"), -- i=2263
      ("00", "1010011001101011", "1101011000101111", "0111110010011010"), -- i=2264
      ("01", "1010011001101011", "1101011000101111", "1101000000111100"), -- i=2265
      ("10", "1010011001101011", "1101011000101111", "1000011000101011"), -- i=2266
      ("11", "1010011001101011", "1101011000101111", "1111011001101111"), -- i=2267
      ("00", "0000101101001100", "0001110010101000", "0010011111110100"), -- i=2268
      ("01", "0000101101001100", "0001110010101000", "1110111010100100"), -- i=2269
      ("10", "0000101101001100", "0001110010101000", "0000100000001000"), -- i=2270
      ("11", "0000101101001100", "0001110010101000", "0001111111101100"), -- i=2271
      ("00", "1101010111111011", "0010110010010100", "0000001010001111"), -- i=2272
      ("01", "1101010111111011", "0010110010010100", "1010100101100111"), -- i=2273
      ("10", "1101010111111011", "0010110010010100", "0000010010010000"), -- i=2274
      ("11", "1101010111111011", "0010110010010100", "1111110111111111"), -- i=2275
      ("00", "0000001111111101", "0100111010101100", "0101001010101001"), -- i=2276
      ("01", "0000001111111101", "0100111010101100", "1011010101010001"), -- i=2277
      ("10", "0000001111111101", "0100111010101100", "0000001010101100"), -- i=2278
      ("11", "0000001111111101", "0100111010101100", "0100111111111101"), -- i=2279
      ("00", "0100001000101000", "0111000011101010", "1011001100010010"), -- i=2280
      ("01", "0100001000101000", "0111000011101010", "1101000100111110"), -- i=2281
      ("10", "0100001000101000", "0111000011101010", "0100000000101000"), -- i=2282
      ("11", "0100001000101000", "0111000011101010", "0111001011101010"), -- i=2283
      ("00", "1011011100011111", "0100101100000001", "0000001000100000"), -- i=2284
      ("01", "1011011100011111", "0100101100000001", "0110110000011110"), -- i=2285
      ("10", "1011011100011111", "0100101100000001", "0000001100000001"), -- i=2286
      ("11", "1011011100011111", "0100101100000001", "1111111100011111"), -- i=2287
      ("00", "0111011001011111", "1110100110000101", "0101111111100100"), -- i=2288
      ("01", "0111011001011111", "1110100110000101", "1000110011011010"), -- i=2289
      ("10", "0111011001011111", "1110100110000101", "0110000000000101"), -- i=2290
      ("11", "0111011001011111", "1110100110000101", "1111111111011111"), -- i=2291
      ("00", "1111101110000011", "0110011000100011", "0110000110100110"), -- i=2292
      ("01", "1111101110000011", "0110011000100011", "1001010101100000"), -- i=2293
      ("10", "1111101110000011", "0110011000100011", "0110001000000011"), -- i=2294
      ("11", "1111101110000011", "0110011000100011", "1111111110100011"), -- i=2295
      ("00", "1110101000110110", "0001010101111010", "1111111110110000"), -- i=2296
      ("01", "1110101000110110", "0001010101111010", "1101010010111100"), -- i=2297
      ("10", "1110101000110110", "0001010101111010", "0000000000110010"), -- i=2298
      ("11", "1110101000110110", "0001010101111010", "1111111101111110"), -- i=2299
      ("00", "1110000010011111", "1001100110000101", "0111101000100100"), -- i=2300
      ("01", "1110000010011111", "1001100110000101", "0100011100011010"), -- i=2301
      ("10", "1110000010011111", "1001100110000101", "1000000010000101"), -- i=2302
      ("11", "1110000010011111", "1001100110000101", "1111100110011111"), -- i=2303
      ("00", "0001110010010100", "1010000101110011", "1011111000000111"), -- i=2304
      ("01", "0001110010010100", "1010000101110011", "0111101100100001"), -- i=2305
      ("10", "0001110010010100", "1010000101110011", "0000000000010000"), -- i=2306
      ("11", "0001110010010100", "1010000101110011", "1011110111110111"), -- i=2307
      ("00", "0100100011001011", "1111000001011110", "0011100100101001"), -- i=2308
      ("01", "0100100011001011", "1111000001011110", "0101100001101101"), -- i=2309
      ("10", "0100100011001011", "1111000001011110", "0100000001001010"), -- i=2310
      ("11", "0100100011001011", "1111000001011110", "1111100011011111"), -- i=2311
      ("00", "0001010001001110", "1100001011001001", "1101011100010111"), -- i=2312
      ("01", "0001010001001110", "1100001011001001", "0101000110000101"), -- i=2313
      ("10", "0001010001001110", "1100001011001001", "0000000001001000"), -- i=2314
      ("11", "0001010001001110", "1100001011001001", "1101011011001111"), -- i=2315
      ("00", "0110010001011111", "0100001010011101", "1010011011111100"), -- i=2316
      ("01", "0110010001011111", "0100001010011101", "0010000111000010"), -- i=2317
      ("10", "0110010001011111", "0100001010011101", "0100000000011101"), -- i=2318
      ("11", "0110010001011111", "0100001010011101", "0110011011011111"), -- i=2319
      ("00", "0111110100111010", "0100100101111100", "1100011010110110"), -- i=2320
      ("01", "0111110100111010", "0100100101111100", "0011001110111110"), -- i=2321
      ("10", "0111110100111010", "0100100101111100", "0100100100111000"), -- i=2322
      ("11", "0111110100111010", "0100100101111100", "0111110101111110"), -- i=2323
      ("00", "0111101000101011", "1100110100101111", "0100011101011010"), -- i=2324
      ("01", "0111101000101011", "1100110100101111", "1010110011111100"), -- i=2325
      ("10", "0111101000101011", "1100110100101111", "0100100000101011"), -- i=2326
      ("11", "0111101000101011", "1100110100101111", "1111111100101111"), -- i=2327
      ("00", "1011110111101100", "1000000011000010", "0011111010101110"), -- i=2328
      ("01", "1011110111101100", "1000000011000010", "0011110100101010"), -- i=2329
      ("10", "1011110111101100", "1000000011000010", "1000000011000000"), -- i=2330
      ("11", "1011110111101100", "1000000011000010", "1011110111101110"), -- i=2331
      ("00", "1010001100111101", "0011000111111011", "1101010100111000"), -- i=2332
      ("01", "1010001100111101", "0011000111111011", "0111000101000010"), -- i=2333
      ("10", "1010001100111101", "0011000111111011", "0010000100111001"), -- i=2334
      ("11", "1010001100111101", "0011000111111011", "1011001111111111"), -- i=2335
      ("00", "1110111110100011", "0110010101000000", "0101010011100011"), -- i=2336
      ("01", "1110111110100011", "0110010101000000", "1000101001100011"), -- i=2337
      ("10", "1110111110100011", "0110010101000000", "0110010100000000"), -- i=2338
      ("11", "1110111110100011", "0110010101000000", "1110111111100011"), -- i=2339
      ("00", "0100000011111011", "1000110101001110", "1100111001001001"), -- i=2340
      ("01", "0100000011111011", "1000110101001110", "1011001110101101"), -- i=2341
      ("10", "0100000011111011", "1000110101001110", "0000000001001010"), -- i=2342
      ("11", "0100000011111011", "1000110101001110", "1100110111111111"), -- i=2343
      ("00", "1001011100010000", "1100111100111010", "0110011001001010"), -- i=2344
      ("01", "1001011100010000", "1100111100111010", "1100011111010110"), -- i=2345
      ("10", "1001011100010000", "1100111100111010", "1000011100010000"), -- i=2346
      ("11", "1001011100010000", "1100111100111010", "1101111100111010"), -- i=2347
      ("00", "1111110111111100", "1001100110001111", "1001011110001011"), -- i=2348
      ("01", "1111110111111100", "1001100110001111", "0110010001101101"), -- i=2349
      ("10", "1111110111111100", "1001100110001111", "1001100110001100"), -- i=2350
      ("11", "1111110111111100", "1001100110001111", "1111110111111111"), -- i=2351
      ("00", "0101101000000010", "1110111000111011", "0100100000111101"), -- i=2352
      ("01", "0101101000000010", "1110111000111011", "0110101111000111"), -- i=2353
      ("10", "0101101000000010", "1110111000111011", "0100101000000010"), -- i=2354
      ("11", "0101101000000010", "1110111000111011", "1111111000111011"), -- i=2355
      ("00", "0001101100101101", "0100110101101110", "0110100010011011"), -- i=2356
      ("01", "0001101100101101", "0100110101101110", "1100110110111111"), -- i=2357
      ("10", "0001101100101101", "0100110101101110", "0000100100101100"), -- i=2358
      ("11", "0001101100101101", "0100110101101110", "0101111101101111"), -- i=2359
      ("00", "1011001100100000", "1101101100001001", "1000111000101001"), -- i=2360
      ("01", "1011001100100000", "1101101100001001", "1101100000010111"), -- i=2361
      ("10", "1011001100100000", "1101101100001001", "1001001100000000"), -- i=2362
      ("11", "1011001100100000", "1101101100001001", "1111101100101001"), -- i=2363
      ("00", "1010010000101000", "1111101111111010", "1010000000100010"), -- i=2364
      ("01", "1010010000101000", "1111101111111010", "1010100000101110"), -- i=2365
      ("10", "1010010000101000", "1111101111111010", "1010000000101000"), -- i=2366
      ("11", "1010010000101000", "1111101111111010", "1111111111111010"), -- i=2367
      ("00", "1101001000111000", "0001001111100000", "1110011000011000"), -- i=2368
      ("01", "1101001000111000", "0001001111100000", "1011111001011000"), -- i=2369
      ("10", "1101001000111000", "0001001111100000", "0001001000100000"), -- i=2370
      ("11", "1101001000111000", "0001001111100000", "1101001111111000"), -- i=2371
      ("00", "1110011011000111", "1100000101000010", "1010100000001001"), -- i=2372
      ("01", "1110011011000111", "1100000101000010", "0010010110000101"), -- i=2373
      ("10", "1110011011000111", "1100000101000010", "1100000001000010"), -- i=2374
      ("11", "1110011011000111", "1100000101000010", "1110011111000111"), -- i=2375
      ("00", "0110110011010111", "0110111001011000", "1101101100101111"), -- i=2376
      ("01", "0110110011010111", "0110111001011000", "1111111001111111"), -- i=2377
      ("10", "0110110011010111", "0110111001011000", "0110110001010000"), -- i=2378
      ("11", "0110110011010111", "0110111001011000", "0110111011011111"), -- i=2379
      ("00", "0011001101011110", "1111000101110000", "0010010011001110"), -- i=2380
      ("01", "0011001101011110", "1111000101110000", "0100000111101110"), -- i=2381
      ("10", "0011001101011110", "1111000101110000", "0011000101010000"), -- i=2382
      ("11", "0011001101011110", "1111000101110000", "1111001101111110"), -- i=2383
      ("00", "0100000000101001", "0110100101011100", "1010100110000101"), -- i=2384
      ("01", "0100000000101001", "0110100101011100", "1101011011001101"), -- i=2385
      ("10", "0100000000101001", "0110100101011100", "0100000000001000"), -- i=2386
      ("11", "0100000000101001", "0110100101011100", "0110100101111101"), -- i=2387
      ("00", "0111110000101011", "0101001110000000", "1100111110101011"), -- i=2388
      ("01", "0111110000101011", "0101001110000000", "0010100010101011"), -- i=2389
      ("10", "0111110000101011", "0101001110000000", "0101000000000000"), -- i=2390
      ("11", "0111110000101011", "0101001110000000", "0111111110101011"), -- i=2391
      ("00", "0110101001001111", "1101000100100100", "0011101101110011"), -- i=2392
      ("01", "0110101001001111", "1101000100100100", "1001100100101011"), -- i=2393
      ("10", "0110101001001111", "1101000100100100", "0100000000000100"), -- i=2394
      ("11", "0110101001001111", "1101000100100100", "1111101101101111"), -- i=2395
      ("00", "1110001111011000", "0010110000001111", "0000111111100111"), -- i=2396
      ("01", "1110001111011000", "0010110000001111", "1011011111001001"), -- i=2397
      ("10", "1110001111011000", "0010110000001111", "0010000000001000"), -- i=2398
      ("11", "1110001111011000", "0010110000001111", "1110111111011111"), -- i=2399
      ("00", "1000111010110100", "0101011000010110", "1110010011001010"), -- i=2400
      ("01", "1000111010110100", "0101011000010110", "0011100010011110"), -- i=2401
      ("10", "1000111010110100", "0101011000010110", "0000011000010100"), -- i=2402
      ("11", "1000111010110100", "0101011000010110", "1101111010110110"), -- i=2403
      ("00", "1010110000110000", "0111111111010000", "0010110000000000"), -- i=2404
      ("01", "1010110000110000", "0111111111010000", "0010110001100000"), -- i=2405
      ("10", "1010110000110000", "0111111111010000", "0010110000010000"), -- i=2406
      ("11", "1010110000110000", "0111111111010000", "1111111111110000"), -- i=2407
      ("00", "1110111000010110", "0000111011110110", "1111110100001100"), -- i=2408
      ("01", "1110111000010110", "0000111011110110", "1101111100100000"), -- i=2409
      ("10", "1110111000010110", "0000111011110110", "0000111000010110"), -- i=2410
      ("11", "1110111000010110", "0000111011110110", "1110111011110110"), -- i=2411
      ("00", "0011111101010100", "1000000010101101", "1100000000000001"), -- i=2412
      ("01", "0011111101010100", "1000000010101101", "1011111010100111"), -- i=2413
      ("10", "0011111101010100", "1000000010101101", "0000000000000100"), -- i=2414
      ("11", "0011111101010100", "1000000010101101", "1011111111111101"), -- i=2415
      ("00", "0011100000110010", "1101110111011101", "0001011000001111"), -- i=2416
      ("01", "0011100000110010", "1101110111011101", "0101101001010101"), -- i=2417
      ("10", "0011100000110010", "1101110111011101", "0001100000010000"), -- i=2418
      ("11", "0011100000110010", "1101110111011101", "1111110111111111"), -- i=2419
      ("00", "0011111100011000", "1100101110101110", "0000101011000110"), -- i=2420
      ("01", "0011111100011000", "1100101110101110", "0111001101101010"), -- i=2421
      ("10", "0011111100011000", "1100101110101110", "0000101100001000"), -- i=2422
      ("11", "0011111100011000", "1100101110101110", "1111111110111110"), -- i=2423
      ("00", "1110001001100000", "0101011011001001", "0011100100101001"), -- i=2424
      ("01", "1110001001100000", "0101011011001001", "1000101110010111"), -- i=2425
      ("10", "1110001001100000", "0101011011001001", "0100001001000000"), -- i=2426
      ("11", "1110001001100000", "0101011011001001", "1111011011101001"), -- i=2427
      ("00", "1001111101010100", "1111100100010010", "1001100001100110"), -- i=2428
      ("01", "1001111101010100", "1111100100010010", "1010011001000010"), -- i=2429
      ("10", "1001111101010100", "1111100100010010", "1001100100010000"), -- i=2430
      ("11", "1001111101010100", "1111100100010010", "1111111101010110"), -- i=2431
      ("00", "0011101110001011", "0001010111001101", "0101000101011000"), -- i=2432
      ("01", "0011101110001011", "0001010111001101", "0010010110111110"), -- i=2433
      ("10", "0011101110001011", "0001010111001101", "0001000110001001"), -- i=2434
      ("11", "0011101110001011", "0001010111001101", "0011111111001111"), -- i=2435
      ("00", "1101000101010010", "0000001101001001", "1101010010011011"), -- i=2436
      ("01", "1101000101010010", "0000001101001001", "1100111000001001"), -- i=2437
      ("10", "1101000101010010", "0000001101001001", "0000000101000000"), -- i=2438
      ("11", "1101000101010010", "0000001101001001", "1101001101011011"), -- i=2439
      ("00", "0100101101000101", "0110101000101100", "1011010101110001"), -- i=2440
      ("01", "0100101101000101", "0110101000101100", "1110000100011001"), -- i=2441
      ("10", "0100101101000101", "0110101000101100", "0100101000000100"), -- i=2442
      ("11", "0100101101000101", "0110101000101100", "0110101101101101"), -- i=2443
      ("00", "1110111110100111", "0011010010110010", "0010010001011001"), -- i=2444
      ("01", "1110111110100111", "0011010010110010", "1011101011110101"), -- i=2445
      ("10", "1110111110100111", "0011010010110010", "0010010010100010"), -- i=2446
      ("11", "1110111110100111", "0011010010110010", "1111111110110111"), -- i=2447
      ("00", "1100011011101010", "1101101011101000", "1010000111010010"), -- i=2448
      ("01", "1100011011101010", "1101101011101000", "1110110000000010"), -- i=2449
      ("10", "1100011011101010", "1101101011101000", "1100001011101000"), -- i=2450
      ("11", "1100011011101010", "1101101011101000", "1101111011101010"), -- i=2451
      ("00", "1010101100010101", "1001111101001110", "0100101001100011"), -- i=2452
      ("01", "1010101100010101", "1001111101001110", "0000101111000111"), -- i=2453
      ("10", "1010101100010101", "1001111101001110", "1000101100000100"), -- i=2454
      ("11", "1010101100010101", "1001111101001110", "1011111101011111"), -- i=2455
      ("00", "0000110100011010", "0101000010010011", "0101110110101101"), -- i=2456
      ("01", "0000110100011010", "0101000010010011", "1011110010000111"), -- i=2457
      ("10", "0000110100011010", "0101000010010011", "0000000000010010"), -- i=2458
      ("11", "0000110100011010", "0101000010010011", "0101110110011011"), -- i=2459
      ("00", "0111001001010001", "1001110011001110", "0000111100011111"), -- i=2460
      ("01", "0111001001010001", "1001110011001110", "1101010110000011"), -- i=2461
      ("10", "0111001001010001", "1001110011001110", "0001000001000000"), -- i=2462
      ("11", "0111001001010001", "1001110011001110", "1111111011011111"), -- i=2463
      ("00", "0010010011110101", "1001111101100010", "1100010001010111"), -- i=2464
      ("01", "0010010011110101", "1001111101100010", "1000010110010011"), -- i=2465
      ("10", "0010010011110101", "1001111101100010", "0000010001100000"), -- i=2466
      ("11", "0010010011110101", "1001111101100010", "1011111111110111"), -- i=2467
      ("00", "1110111111001000", "0111100010100110", "0110100001101110"), -- i=2468
      ("01", "1110111111001000", "0111100010100110", "0111011100100010"), -- i=2469
      ("10", "1110111111001000", "0111100010100110", "0110100010000000"), -- i=2470
      ("11", "1110111111001000", "0111100010100110", "1111111111101110"), -- i=2471
      ("00", "0011001111011011", "1100001111011101", "1111011110111000"), -- i=2472
      ("01", "0011001111011011", "1100001111011101", "0110111111111110"), -- i=2473
      ("10", "0011001111011011", "1100001111011101", "0000001111011001"), -- i=2474
      ("11", "0011001111011011", "1100001111011101", "1111001111011111"), -- i=2475
      ("00", "1000000110111100", "0011000100010011", "1011001011001111"), -- i=2476
      ("01", "1000000110111100", "0011000100010011", "0101000010101001"), -- i=2477
      ("10", "1000000110111100", "0011000100010011", "0000000100010000"), -- i=2478
      ("11", "1000000110111100", "0011000100010011", "1011000110111111"), -- i=2479
      ("00", "1011100110100110", "0110001110100001", "0001110101000111"), -- i=2480
      ("01", "1011100110100110", "0110001110100001", "0101011000000101"), -- i=2481
      ("10", "1011100110100110", "0110001110100001", "0010000110100000"), -- i=2482
      ("11", "1011100110100110", "0110001110100001", "1111101110100111"), -- i=2483
      ("00", "1100001001001001", "0010111100110011", "1111000101111100"), -- i=2484
      ("01", "1100001001001001", "0010111100110011", "1001001100010110"), -- i=2485
      ("10", "1100001001001001", "0010111100110011", "0000001000000001"), -- i=2486
      ("11", "1100001001001001", "0010111100110011", "1110111101111011"), -- i=2487
      ("00", "0010100010100011", "0000101100010000", "0011001110110011"), -- i=2488
      ("01", "0010100010100011", "0000101100010000", "0001110110010011"), -- i=2489
      ("10", "0010100010100011", "0000101100010000", "0000100000000000"), -- i=2490
      ("11", "0010100010100011", "0000101100010000", "0010101110110011"), -- i=2491
      ("00", "1000111001000111", "1111000110101001", "0111111111110000"), -- i=2492
      ("01", "1000111001000111", "1111000110101001", "1001110010011110"), -- i=2493
      ("10", "1000111001000111", "1111000110101001", "1000000000000001"), -- i=2494
      ("11", "1000111001000111", "1111000110101001", "1111111111101111"), -- i=2495
      ("00", "0001101110101111", "0010111111110000", "0100101110011111"), -- i=2496
      ("01", "0001101110101111", "0010111111110000", "1110101110111111"), -- i=2497
      ("10", "0001101110101111", "0010111111110000", "0000101110100000"), -- i=2498
      ("11", "0001101110101111", "0010111111110000", "0011111111111111"), -- i=2499
      ("00", "0011101011111110", "1110100001101111", "0010001101101101"), -- i=2500
      ("01", "0011101011111110", "1110100001101111", "0101001010001111"), -- i=2501
      ("10", "0011101011111110", "1110100001101111", "0010100001101110"), -- i=2502
      ("11", "0011101011111110", "1110100001101111", "1111101011111111"), -- i=2503
      ("00", "1000001001000111", "0011100001000101", "1011101010001100"), -- i=2504
      ("01", "1000001001000111", "0011100001000101", "0100101000000010"), -- i=2505
      ("10", "1000001001000111", "0011100001000101", "0000000001000101"), -- i=2506
      ("11", "1000001001000111", "0011100001000101", "1011101001000111"), -- i=2507
      ("00", "1101010000100110", "0010101110110110", "1111111111011100"), -- i=2508
      ("01", "1101010000100110", "0010101110110110", "1010100001110000"), -- i=2509
      ("10", "1101010000100110", "0010101110110110", "0000000000100110"), -- i=2510
      ("11", "1101010000100110", "0010101110110110", "1111111110110110"), -- i=2511
      ("00", "1001011101111001", "1010001111101011", "0011101101100100"), -- i=2512
      ("01", "1001011101111001", "1010001111101011", "1111001110001110"), -- i=2513
      ("10", "1001011101111001", "1010001111101011", "1000001101101001"), -- i=2514
      ("11", "1001011101111001", "1010001111101011", "1011011111111011"), -- i=2515
      ("00", "0100110010111101", "0100101100010100", "1001011111010001"), -- i=2516
      ("01", "0100110010111101", "0100101100010100", "0000000110101001"), -- i=2517
      ("10", "0100110010111101", "0100101100010100", "0100100000010100"), -- i=2518
      ("11", "0100110010111101", "0100101100010100", "0100111110111101"), -- i=2519
      ("00", "0101110111110100", "1111111011001010", "0101110010111110"), -- i=2520
      ("01", "0101110111110100", "1111111011001010", "0101111100101010"), -- i=2521
      ("10", "0101110111110100", "1111111011001010", "0101110011000000"), -- i=2522
      ("11", "0101110111110100", "1111111011001010", "1111111111111110"), -- i=2523
      ("00", "1000011010001111", "0010110101010100", "1011001111100011"), -- i=2524
      ("01", "1000011010001111", "0010110101010100", "0101100100111011"), -- i=2525
      ("10", "1000011010001111", "0010110101010100", "0000010000000100"), -- i=2526
      ("11", "1000011010001111", "0010110101010100", "1010111111011111"), -- i=2527
      ("00", "1010100010110001", "0111000010010111", "0001100101001000"), -- i=2528
      ("01", "1010100010110001", "0111000010010111", "0011100000011010"), -- i=2529
      ("10", "1010100010110001", "0111000010010111", "0010000010010001"), -- i=2530
      ("11", "1010100010110001", "0111000010010111", "1111100010110111"), -- i=2531
      ("00", "1111010110001101", "1101110010100100", "1101001000110001"), -- i=2532
      ("01", "1111010110001101", "1101110010100100", "0001100011101001"), -- i=2533
      ("10", "1111010110001101", "1101110010100100", "1101010010000100"), -- i=2534
      ("11", "1111010110001101", "1101110010100100", "1111110110101101"), -- i=2535
      ("00", "0110110011101101", "1001011001111110", "0000001101101011"), -- i=2536
      ("01", "0110110011101101", "1001011001111110", "1101011001101111"), -- i=2537
      ("10", "0110110011101101", "1001011001111110", "0000010001101100"), -- i=2538
      ("11", "0110110011101101", "1001011001111110", "1111111011111111"), -- i=2539
      ("00", "0110110101000111", "0010010111111110", "1001001101000101"), -- i=2540
      ("01", "0110110101000111", "0010010111111110", "0100011101001001"), -- i=2541
      ("10", "0110110101000111", "0010010111111110", "0010010101000110"), -- i=2542
      ("11", "0110110101000111", "0010010111111110", "0110110111111111"), -- i=2543
      ("00", "0011011101101111", "1101001000110110", "0000100110100101"), -- i=2544
      ("01", "0011011101101111", "1101001000110110", "0110010100111001"), -- i=2545
      ("10", "0011011101101111", "1101001000110110", "0001001000100110"), -- i=2546
      ("11", "0011011101101111", "1101001000110110", "1111011101111111"), -- i=2547
      ("00", "0101100000110010", "0010010111110111", "0111111000101001"), -- i=2548
      ("01", "0101100000110010", "0010010111110111", "0011001000111011"), -- i=2549
      ("10", "0101100000110010", "0010010111110111", "0000000000110010"), -- i=2550
      ("11", "0101100000110010", "0010010111110111", "0111110111110111"), -- i=2551
      ("00", "0010010001010111", "0110000101010010", "1000010110101001"), -- i=2552
      ("01", "0010010001010111", "0110000101010010", "1100001100000101"), -- i=2553
      ("10", "0010010001010111", "0110000101010010", "0010000001010010"), -- i=2554
      ("11", "0010010001010111", "0110000101010010", "0110010101010111"), -- i=2555
      ("00", "0011000101111010", "0011100001101110", "0110100111101000"), -- i=2556
      ("01", "0011000101111010", "0011100001101110", "1111100100001100"), -- i=2557
      ("10", "0011000101111010", "0011100001101110", "0011000001101010"), -- i=2558
      ("11", "0011000101111010", "0011100001101110", "0011100101111110"), -- i=2559
      ("00", "1010010111101010", "0101111011001000", "0000010010110010"), -- i=2560
      ("01", "1010010111101010", "0101111011001000", "0100011100100010"), -- i=2561
      ("10", "1010010111101010", "0101111011001000", "0000010011001000"), -- i=2562
      ("11", "1010010111101010", "0101111011001000", "1111111111101010"), -- i=2563
      ("00", "1001101110010110", "0100001110101011", "1101111101000001"), -- i=2564
      ("01", "1001101110010110", "0100001110101011", "0101011111101011"), -- i=2565
      ("10", "1001101110010110", "0100001110101011", "0000001110000010"), -- i=2566
      ("11", "1001101110010110", "0100001110101011", "1101101110111111"), -- i=2567
      ("00", "1011110000011011", "0100100000001111", "0000010000101010"), -- i=2568
      ("01", "1011110000011011", "0100100000001111", "0111010000001100"), -- i=2569
      ("10", "1011110000011011", "0100100000001111", "0000100000001011"), -- i=2570
      ("11", "1011110000011011", "0100100000001111", "1111110000011111"), -- i=2571
      ("00", "1101011011101000", "0000001011110010", "1101100111011010"), -- i=2572
      ("01", "1101011011101000", "0000001011110010", "1101001111110110"), -- i=2573
      ("10", "1101011011101000", "0000001011110010", "0000001011100000"), -- i=2574
      ("11", "1101011011101000", "0000001011110010", "1101011011111010"), -- i=2575
      ("00", "1111101111000111", "1011111001000111", "1011101000001110"), -- i=2576
      ("01", "1111101111000111", "1011111001000111", "0011110110000000"), -- i=2577
      ("10", "1111101111000111", "1011111001000111", "1011101001000111"), -- i=2578
      ("11", "1111101111000111", "1011111001000111", "1111111111000111"), -- i=2579
      ("00", "1010110011111111", "1100011110011011", "0111010010011010"), -- i=2580
      ("01", "1010110011111111", "1100011110011011", "1110010101100100"), -- i=2581
      ("10", "1010110011111111", "1100011110011011", "1000010010011011"), -- i=2582
      ("11", "1010110011111111", "1100011110011011", "1110111111111111"), -- i=2583
      ("00", "1110100111011111", "0000001101000110", "1110110100100101"), -- i=2584
      ("01", "1110100111011111", "0000001101000110", "1110011010011001"), -- i=2585
      ("10", "1110100111011111", "0000001101000110", "0000000101000110"), -- i=2586
      ("11", "1110100111011111", "0000001101000110", "1110101111011111"), -- i=2587
      ("00", "0001111001101011", "0010001100110010", "0100000110011101"), -- i=2588
      ("01", "0001111001101011", "0010001100110010", "1111101100111001"), -- i=2589
      ("10", "0001111001101011", "0010001100110010", "0000001000100010"), -- i=2590
      ("11", "0001111001101011", "0010001100110010", "0011111101111011"), -- i=2591
      ("00", "1011101111111001", "0010000110001111", "1101110110001000"), -- i=2592
      ("01", "1011101111111001", "0010000110001111", "1001101001101010"), -- i=2593
      ("10", "1011101111111001", "0010000110001111", "0010000110001001"), -- i=2594
      ("11", "1011101111111001", "0010000110001111", "1011101111111111"), -- i=2595
      ("00", "0100001000011101", "0001000000110111", "0101001001010100"), -- i=2596
      ("01", "0100001000011101", "0001000000110111", "0011000111100110"), -- i=2597
      ("10", "0100001000011101", "0001000000110111", "0000000000010101"), -- i=2598
      ("11", "0100001000011101", "0001000000110111", "0101001000111111"), -- i=2599
      ("00", "1000010100001001", "1100010101110101", "0100101001111110"), -- i=2600
      ("01", "1000010100001001", "1100010101110101", "1011111110010100"), -- i=2601
      ("10", "1000010100001001", "1100010101110101", "1000010100000001"), -- i=2602
      ("11", "1000010100001001", "1100010101110101", "1100010101111101"), -- i=2603
      ("00", "1100111011001110", "0111101001101011", "0100100100111001"), -- i=2604
      ("01", "1100111011001110", "0111101001101011", "0101010001100011"), -- i=2605
      ("10", "1100111011001110", "0111101001101011", "0100101001001010"), -- i=2606
      ("11", "1100111011001110", "0111101001101011", "1111111011101111"), -- i=2607
      ("00", "0011001000110000", "1000110100000010", "1011111100110010"), -- i=2608
      ("01", "0011001000110000", "1000110100000010", "1010010100101110"), -- i=2609
      ("10", "0011001000110000", "1000110100000010", "0000000000000000"), -- i=2610
      ("11", "0011001000110000", "1000110100000010", "1011111100110010"), -- i=2611
      ("00", "1011011111101011", "0111101011100000", "0011001011001011"), -- i=2612
      ("01", "1011011111101011", "0111101011100000", "0011110100001011"), -- i=2613
      ("10", "1011011111101011", "0111101011100000", "0011001011100000"), -- i=2614
      ("11", "1011011111101011", "0111101011100000", "1111111111101011"), -- i=2615
      ("00", "1000000011100011", "1111101101100010", "0111110001000101"), -- i=2616
      ("01", "1000000011100011", "1111101101100010", "1000010110000001"), -- i=2617
      ("10", "1000000011100011", "1111101101100010", "1000000001100010"), -- i=2618
      ("11", "1000000011100011", "1111101101100010", "1111101111100011"), -- i=2619
      ("00", "0010000011110100", "0011011100100001", "0101100000010101"), -- i=2620
      ("01", "0010000011110100", "0011011100100001", "1110100111010011"), -- i=2621
      ("10", "0010000011110100", "0011011100100001", "0010000000100000"), -- i=2622
      ("11", "0010000011110100", "0011011100100001", "0011011111110101"), -- i=2623
      ("00", "0100010011100110", "0100101111011011", "1001000011000001"), -- i=2624
      ("01", "0100010011100110", "0100101111011011", "1111100100001011"), -- i=2625
      ("10", "0100010011100110", "0100101111011011", "0100000011000010"), -- i=2626
      ("11", "0100010011100110", "0100101111011011", "0100111111111111"), -- i=2627
      ("00", "1010101101100001", "0001011000110001", "1100000110010010"), -- i=2628
      ("01", "1010101101100001", "0001011000110001", "1001010100110000"), -- i=2629
      ("10", "1010101101100001", "0001011000110001", "0000001000100001"), -- i=2630
      ("11", "1010101101100001", "0001011000110001", "1011111101110001"), -- i=2631
      ("00", "1110100111001100", "0001011110101001", "0000000101110101"), -- i=2632
      ("01", "1110100111001100", "0001011110101001", "1101001000100011"), -- i=2633
      ("10", "1110100111001100", "0001011110101001", "0000000110001000"), -- i=2634
      ("11", "1110100111001100", "0001011110101001", "1111111111101101"), -- i=2635
      ("00", "1100110001011100", "1110100100111101", "1011010110011001"), -- i=2636
      ("01", "1100110001011100", "1110100100111101", "1110001100011111"), -- i=2637
      ("10", "1100110001011100", "1110100100111101", "1100100000011100"), -- i=2638
      ("11", "1100110001011100", "1110100100111101", "1110110101111101"), -- i=2639
      ("00", "0001100011111100", "0010000100110101", "0011101000110001"), -- i=2640
      ("01", "0001100011111100", "0010000100110101", "1111011111000111"), -- i=2641
      ("10", "0001100011111100", "0010000100110101", "0000000000110100"), -- i=2642
      ("11", "0001100011111100", "0010000100110101", "0011100111111101"), -- i=2643
      ("00", "0110100100000010", "1011100100110110", "0010001000111000"), -- i=2644
      ("01", "0110100100000010", "1011100100110110", "1010111111001100"), -- i=2645
      ("10", "0110100100000010", "1011100100110110", "0010100100000010"), -- i=2646
      ("11", "0110100100000010", "1011100100110110", "1111100100110110"), -- i=2647
      ("00", "1101001001111010", "1001111010000001", "0111000011111011"), -- i=2648
      ("01", "1101001001111010", "1001111010000001", "0011001111111001"), -- i=2649
      ("10", "1101001001111010", "1001111010000001", "1001001000000000"), -- i=2650
      ("11", "1101001001111010", "1001111010000001", "1101111011111011"), -- i=2651
      ("00", "0111000011101110", "0010010110101011", "1001011010011001"), -- i=2652
      ("01", "0111000011101110", "0010010110101011", "0100101101000011"), -- i=2653
      ("10", "0111000011101110", "0010010110101011", "0010000010101010"), -- i=2654
      ("11", "0111000011101110", "0010010110101011", "0111010111101111"), -- i=2655
      ("00", "0001001111100001", "0000101111001011", "0001111110101100"), -- i=2656
      ("01", "0001001111100001", "0000101111001011", "0000100000010110"), -- i=2657
      ("10", "0001001111100001", "0000101111001011", "0000001111000001"), -- i=2658
      ("11", "0001001111100001", "0000101111001011", "0001101111101011"), -- i=2659
      ("00", "1001000000110100", "1010010010100110", "0011010011011010"), -- i=2660
      ("01", "1001000000110100", "1010010010100110", "1110101110001110"), -- i=2661
      ("10", "1001000000110100", "1010010010100110", "1000000000100100"), -- i=2662
      ("11", "1001000000110100", "1010010010100110", "1011010010110110"), -- i=2663
      ("00", "0101111001010111", "1110011010101111", "0100010100000110"), -- i=2664
      ("01", "0101111001010111", "1110011010101111", "0111011110101000"), -- i=2665
      ("10", "0101111001010111", "1110011010101111", "0100011000000111"), -- i=2666
      ("11", "0101111001010111", "1110011010101111", "1111111011111111"), -- i=2667
      ("00", "0101101100100110", "0111111001011111", "1101100110000101"), -- i=2668
      ("01", "0101101100100110", "0111111001011111", "1101110011000111"), -- i=2669
      ("10", "0101101100100110", "0111111001011111", "0101101000000110"), -- i=2670
      ("11", "0101101100100110", "0111111001011111", "0111111101111111"), -- i=2671
      ("00", "0000100101100010", "1011000101100010", "1011101011000100"), -- i=2672
      ("01", "0000100101100010", "1011000101100010", "0101100000000000"), -- i=2673
      ("10", "0000100101100010", "1011000101100010", "0000000101100010"), -- i=2674
      ("11", "0000100101100010", "1011000101100010", "1011100101100010"), -- i=2675
      ("00", "1000011101110101", "0001001100000000", "1001101001110101"), -- i=2676
      ("01", "1000011101110101", "0001001100000000", "0111010001110101"), -- i=2677
      ("10", "1000011101110101", "0001001100000000", "0000001100000000"), -- i=2678
      ("11", "1000011101110101", "0001001100000000", "1001011101110101"), -- i=2679
      ("00", "0101010111101111", "0100010010110010", "1001101010100001"), -- i=2680
      ("01", "0101010111101111", "0100010010110010", "0001000100111101"), -- i=2681
      ("10", "0101010111101111", "0100010010110010", "0100010010100010"), -- i=2682
      ("11", "0101010111101111", "0100010010110010", "0101010111111111"), -- i=2683
      ("00", "1101111110010000", "1101001111011001", "1011001101101001"), -- i=2684
      ("01", "1101111110010000", "1101001111011001", "0000101110110111"), -- i=2685
      ("10", "1101111110010000", "1101001111011001", "1101001110010000"), -- i=2686
      ("11", "1101111110010000", "1101001111011001", "1101111111011001"), -- i=2687
      ("00", "1010000111110110", "1100011011110101", "0110100011101011"), -- i=2688
      ("01", "1010000111110110", "1100011011110101", "1101101100000001"), -- i=2689
      ("10", "1010000111110110", "1100011011110101", "1000000011110100"), -- i=2690
      ("11", "1010000111110110", "1100011011110101", "1110011111110111"), -- i=2691
      ("00", "1001111001011100", "0101110010101101", "1111101100001001"), -- i=2692
      ("01", "1001111001011100", "0101110010101101", "0100000110101111"), -- i=2693
      ("10", "1001111001011100", "0101110010101101", "0001110000001100"), -- i=2694
      ("11", "1001111001011100", "0101110010101101", "1101111011111101"), -- i=2695
      ("00", "1111001001110001", "1001010100011110", "1000011110001111"), -- i=2696
      ("01", "1111001001110001", "1001010100011110", "0101110101010011"), -- i=2697
      ("10", "1111001001110001", "1001010100011110", "1001000000010000"), -- i=2698
      ("11", "1111001001110001", "1001010100011110", "1111011101111111"), -- i=2699
      ("00", "1100101010010010", "0100010100010101", "0000111110100111"), -- i=2700
      ("01", "1100101010010010", "0100010100010101", "1000010101111101"), -- i=2701
      ("10", "1100101010010010", "0100010100010101", "0100000000010000"), -- i=2702
      ("11", "1100101010010010", "0100010100010101", "1100111110010111"), -- i=2703
      ("00", "0100011010110010", "0000101010000111", "0101000100111001"), -- i=2704
      ("01", "0100011010110010", "0000101010000111", "0011110000101011"), -- i=2705
      ("10", "0100011010110010", "0000101010000111", "0000001010000010"), -- i=2706
      ("11", "0100011010110010", "0000101010000111", "0100111010110111"), -- i=2707
      ("00", "1111101001110011", "1001010100000101", "1000111101111000"), -- i=2708
      ("01", "1111101001110011", "1001010100000101", "0110010101101110"), -- i=2709
      ("10", "1111101001110011", "1001010100000101", "1001000000000001"), -- i=2710
      ("11", "1111101001110011", "1001010100000101", "1111111101110111"), -- i=2711
      ("00", "1100110101000010", "0101101100110110", "0010100001111000"), -- i=2712
      ("01", "1100110101000010", "0101101100110110", "0111001000001100"), -- i=2713
      ("10", "1100110101000010", "0101101100110110", "0100100100000010"), -- i=2714
      ("11", "1100110101000010", "0101101100110110", "1101111101110110"), -- i=2715
      ("00", "1010000110010001", "0100001011110110", "1110010010000111"), -- i=2716
      ("01", "1010000110010001", "0100001011110110", "0101111010011011"), -- i=2717
      ("10", "1010000110010001", "0100001011110110", "0000000010010000"), -- i=2718
      ("11", "1010000110010001", "0100001011110110", "1110001111110111"), -- i=2719
      ("00", "0001111111000111", "1010001110110011", "1100001101111010"), -- i=2720
      ("01", "0001111111000111", "1010001110110011", "0111110000010100"), -- i=2721
      ("10", "0001111111000111", "1010001110110011", "0000001110000011"), -- i=2722
      ("11", "0001111111000111", "1010001110110011", "1011111111110111"), -- i=2723
      ("00", "1010101111100100", "1100010101010101", "0111000100111001"), -- i=2724
      ("01", "1010101111100100", "1100010101010101", "1110011010001111"), -- i=2725
      ("10", "1010101111100100", "1100010101010101", "1000000101000100"), -- i=2726
      ("11", "1010101111100100", "1100010101010101", "1110111111110101"), -- i=2727
      ("00", "0010000010101110", "1110100010101001", "0000100101010111"), -- i=2728
      ("01", "0010000010101110", "1110100010101001", "0011100000000101"), -- i=2729
      ("10", "0010000010101110", "1110100010101001", "0010000010101000"), -- i=2730
      ("11", "0010000010101110", "1110100010101001", "1110100010101111"), -- i=2731
      ("00", "1011001001101010", "1000110000011110", "0011111010001000"), -- i=2732
      ("01", "1011001001101010", "1000110000011110", "0010011001001100"), -- i=2733
      ("10", "1011001001101010", "1000110000011110", "1000000000001010"), -- i=2734
      ("11", "1011001001101010", "1000110000011110", "1011111001111110"), -- i=2735
      ("00", "1111001010010100", "1111111111101010", "1111001001111110"), -- i=2736
      ("01", "1111001010010100", "1111111111101010", "1111001010101010"), -- i=2737
      ("10", "1111001010010100", "1111111111101010", "1111001010000000"), -- i=2738
      ("11", "1111001010010100", "1111111111101010", "1111111111111110"), -- i=2739
      ("00", "1000011011111101", "0010101011010100", "1011000111010001"), -- i=2740
      ("01", "1000011011111101", "0010101011010100", "0101110000101001"), -- i=2741
      ("10", "1000011011111101", "0010101011010100", "0000001011010100"), -- i=2742
      ("11", "1000011011111101", "0010101011010100", "1010111011111101"), -- i=2743
      ("00", "1100011010011110", "0100001110010100", "0000101000110010"), -- i=2744
      ("01", "1100011010011110", "0100001110010100", "1000001100001010"), -- i=2745
      ("10", "1100011010011110", "0100001110010100", "0100001010010100"), -- i=2746
      ("11", "1100011010011110", "0100001110010100", "1100011110011110"), -- i=2747
      ("00", "0010111000111001", "0001011000111101", "0100010001110110"), -- i=2748
      ("01", "0010111000111001", "0001011000111101", "0001011111111100"), -- i=2749
      ("10", "0010111000111001", "0001011000111101", "0000011000111001"), -- i=2750
      ("11", "0010111000111001", "0001011000111101", "0011111000111101"), -- i=2751
      ("00", "1110110001001101", "0111111101101010", "0110101110110111"), -- i=2752
      ("01", "1110110001001101", "0111111101101010", "0110110011100011"), -- i=2753
      ("10", "1110110001001101", "0111111101101010", "0110110001001000"), -- i=2754
      ("11", "1110110001001101", "0111111101101010", "1111111101101111"), -- i=2755
      ("00", "1001111101111111", "0001110010001010", "1011110000001001"), -- i=2756
      ("01", "1001111101111111", "0001110010001010", "1000001011110101"), -- i=2757
      ("10", "1001111101111111", "0001110010001010", "0001110000001010"), -- i=2758
      ("11", "1001111101111111", "0001110010001010", "1001111111111111"), -- i=2759
      ("00", "1010001001101110", "1011111110101011", "0110001000011001"), -- i=2760
      ("01", "1010001001101110", "1011111110101011", "1110001011000011"), -- i=2761
      ("10", "1010001001101110", "1011111110101011", "1010001000101010"), -- i=2762
      ("11", "1010001001101110", "1011111110101011", "1011111111101111"), -- i=2763
      ("00", "1100110001111100", "0010100111011000", "1111011001010100"), -- i=2764
      ("01", "1100110001111100", "0010100111011000", "1010001010100100"), -- i=2765
      ("10", "1100110001111100", "0010100111011000", "0000100001011000"), -- i=2766
      ("11", "1100110001111100", "0010100111011000", "1110110111111100"), -- i=2767
      ("00", "1010011000111100", "1000011111100100", "0010111000100000"), -- i=2768
      ("01", "1010011000111100", "1000011111100100", "0001111001011000"), -- i=2769
      ("10", "1010011000111100", "1000011111100100", "1000011000100100"), -- i=2770
      ("11", "1010011000111100", "1000011111100100", "1010011111111100"), -- i=2771
      ("00", "1000001011001010", "0111111000110001", "0000000011111011"), -- i=2772
      ("01", "1000001011001010", "0111111000110001", "0000010010011001"), -- i=2773
      ("10", "1000001011001010", "0111111000110001", "0000001000000000"), -- i=2774
      ("11", "1000001011001010", "0111111000110001", "1111111011111011"), -- i=2775
      ("00", "0110001011010011", "0111111110011101", "1110001001110000"), -- i=2776
      ("01", "0110001011010011", "0111111110011101", "1110001100110110"), -- i=2777
      ("10", "0110001011010011", "0111111110011101", "0110001010010001"), -- i=2778
      ("11", "0110001011010011", "0111111110011101", "0111111111011111"), -- i=2779
      ("00", "1011001110000010", "0011010101111101", "1110100011111111"), -- i=2780
      ("01", "1011001110000010", "0011010101111101", "0111111000000101"), -- i=2781
      ("10", "1011001110000010", "0011010101111101", "0011000100000000"), -- i=2782
      ("11", "1011001110000010", "0011010101111101", "1011011111111111"), -- i=2783
      ("00", "1111000010001010", "1101000111011000", "1100001001100010"), -- i=2784
      ("01", "1111000010001010", "1101000111011000", "0001111010110010"), -- i=2785
      ("10", "1111000010001010", "1101000111011000", "1101000010001000"), -- i=2786
      ("11", "1111000010001010", "1101000111011000", "1111000111011010"), -- i=2787
      ("00", "1000110111011010", "1110010100000011", "0111001011011101"), -- i=2788
      ("01", "1000110111011010", "1110010100000011", "1010100011010111"), -- i=2789
      ("10", "1000110111011010", "1110010100000011", "1000010100000010"), -- i=2790
      ("11", "1000110111011010", "1110010100000011", "1110110111011011"), -- i=2791
      ("00", "1100100011010010", "0101001110101110", "0001110010000000"), -- i=2792
      ("01", "1100100011010010", "0101001110101110", "0111010100100100"), -- i=2793
      ("10", "1100100011010010", "0101001110101110", "0100000010000010"), -- i=2794
      ("11", "1100100011010010", "0101001110101110", "1101101111111110"), -- i=2795
      ("00", "1010001100110011", "0001110101110000", "1100000010100011"), -- i=2796
      ("01", "1010001100110011", "0001110101110000", "1000010111000011"), -- i=2797
      ("10", "1010001100110011", "0001110101110000", "0000000100110000"), -- i=2798
      ("11", "1010001100110011", "0001110101110000", "1011111101110011"), -- i=2799
      ("00", "0011000010101001", "0000010110100111", "0011011001010000"), -- i=2800
      ("01", "0011000010101001", "0000010110100111", "0010101100000010"), -- i=2801
      ("10", "0011000010101001", "0000010110100111", "0000000010100001"), -- i=2802
      ("11", "0011000010101001", "0000010110100111", "0011010110101111"), -- i=2803
      ("00", "1111110000011000", "1101001110000001", "1100111110011001"), -- i=2804
      ("01", "1111110000011000", "1101001110000001", "0010100010010111"), -- i=2805
      ("10", "1111110000011000", "1101001110000001", "1101000000000000"), -- i=2806
      ("11", "1111110000011000", "1101001110000001", "1111111110011001"), -- i=2807
      ("00", "1110000011010001", "1010101001111010", "1000101101001011"), -- i=2808
      ("01", "1110000011010001", "1010101001111010", "0011011001010111"), -- i=2809
      ("10", "1110000011010001", "1010101001111010", "1010000001010000"), -- i=2810
      ("11", "1110000011010001", "1010101001111010", "1110101011111011"), -- i=2811
      ("00", "1001111100101100", "0000110011001001", "1010101111110101"), -- i=2812
      ("01", "1001111100101100", "0000110011001001", "1001001001100011"), -- i=2813
      ("10", "1001111100101100", "0000110011001001", "0000110000001000"), -- i=2814
      ("11", "1001111100101100", "0000110011001001", "1001111111101101"), -- i=2815
      ("00", "0110000001001000", "1111110101010111", "0101110110011111"), -- i=2816
      ("01", "0110000001001000", "1111110101010111", "0110001011110001"), -- i=2817
      ("10", "0110000001001000", "1111110101010111", "0110000001000000"), -- i=2818
      ("11", "0110000001001000", "1111110101010111", "1111110101011111"), -- i=2819
      ("00", "1000101111111100", "1011000100101100", "0011110100101000"), -- i=2820
      ("01", "1000101111111100", "1011000100101100", "1101101011010000"), -- i=2821
      ("10", "1000101111111100", "1011000100101100", "1000000100101100"), -- i=2822
      ("11", "1000101111111100", "1011000100101100", "1011101111111100"), -- i=2823
      ("00", "1101101010111000", "1000100011111001", "0110001110110001"), -- i=2824
      ("01", "1101101010111000", "1000100011111001", "0101000110111111"), -- i=2825
      ("10", "1101101010111000", "1000100011111001", "1000100010111000"), -- i=2826
      ("11", "1101101010111000", "1000100011111001", "1101101011111001"), -- i=2827
      ("00", "1001010100101101", "0000110100001000", "1010001000110101"), -- i=2828
      ("01", "1001010100101101", "0000110100001000", "1000100000100101"), -- i=2829
      ("10", "1001010100101101", "0000110100001000", "0000010100001000"), -- i=2830
      ("11", "1001010100101101", "0000110100001000", "1001110100101101"), -- i=2831
      ("00", "1111100111011111", "0100000000001011", "0011100111101010"), -- i=2832
      ("01", "1111100111011111", "0100000000001011", "1011100111010100"), -- i=2833
      ("10", "1111100111011111", "0100000000001011", "0100000000001011"), -- i=2834
      ("11", "1111100111011111", "0100000000001011", "1111100111011111"), -- i=2835
      ("00", "1101011010001010", "0110001100110000", "0011100110111010"), -- i=2836
      ("01", "1101011010001010", "0110001100110000", "0111001101011010"), -- i=2837
      ("10", "1101011010001010", "0110001100110000", "0100001000000000"), -- i=2838
      ("11", "1101011010001010", "0110001100110000", "1111011110111010"), -- i=2839
      ("00", "0110111000100011", "1011111010110000", "0010110011010011"), -- i=2840
      ("01", "0110111000100011", "1011111010110000", "1010111101110011"), -- i=2841
      ("10", "0110111000100011", "1011111010110000", "0010111000100000"), -- i=2842
      ("11", "0110111000100011", "1011111010110000", "1111111010110011"), -- i=2843
      ("00", "1011110011011100", "1110100100011101", "1010010111111001"), -- i=2844
      ("01", "1011110011011100", "1110100100011101", "1101001110111111"), -- i=2845
      ("10", "1011110011011100", "1110100100011101", "1010100000011100"), -- i=2846
      ("11", "1011110011011100", "1110100100011101", "1111110111011101"), -- i=2847
      ("00", "0101111111010000", "1000110000101111", "1110101111111111"), -- i=2848
      ("01", "0101111111010000", "1000110000101111", "1101001110100001"), -- i=2849
      ("10", "0101111111010000", "1000110000101111", "0000110000000000"), -- i=2850
      ("11", "0101111111010000", "1000110000101111", "1101111111111111"), -- i=2851
      ("00", "1011011010011100", "1010101100001011", "0110000110100111"), -- i=2852
      ("01", "1011011010011100", "1010101100001011", "0000101110010001"), -- i=2853
      ("10", "1011011010011100", "1010101100001011", "1010001000001000"), -- i=2854
      ("11", "1011011010011100", "1010101100001011", "1011111110011111"), -- i=2855
      ("00", "1111011110110011", "1100101100010111", "1100001011001010"), -- i=2856
      ("01", "1111011110110011", "1100101100010111", "0010110010011100"), -- i=2857
      ("10", "1111011110110011", "1100101100010111", "1100001100010011"), -- i=2858
      ("11", "1111011110110011", "1100101100010111", "1111111110110111"), -- i=2859
      ("00", "1010110111011011", "0010000011100010", "1100111010111101"), -- i=2860
      ("01", "1010110111011011", "0010000011100010", "1000110011111001"), -- i=2861
      ("10", "1010110111011011", "0010000011100010", "0010000011000010"), -- i=2862
      ("11", "1010110111011011", "0010000011100010", "1010110111111011"), -- i=2863
      ("00", "1000101100011011", "1000010101011010", "0001000001110101"), -- i=2864
      ("01", "1000101100011011", "1000010101011010", "0000010111000001"), -- i=2865
      ("10", "1000101100011011", "1000010101011010", "1000000100011010"), -- i=2866
      ("11", "1000101100011011", "1000010101011010", "1000111101011011"), -- i=2867
      ("00", "0101110100000011", "1011000000011100", "0000110100011111"), -- i=2868
      ("01", "0101110100000011", "1011000000011100", "1010110011100111"), -- i=2869
      ("10", "0101110100000011", "1011000000011100", "0001000000000000"), -- i=2870
      ("11", "0101110100000011", "1011000000011100", "1111110100011111"), -- i=2871
      ("00", "1011110001100111", "0010100100110011", "1110010110011010"), -- i=2872
      ("01", "1011110001100111", "0010100100110011", "1001001100110100"), -- i=2873
      ("10", "1011110001100111", "0010100100110011", "0010100000100011"), -- i=2874
      ("11", "1011110001100111", "0010100100110011", "1011110101110111"), -- i=2875
      ("00", "0110100100110101", "1111001000001100", "0101101101000001"), -- i=2876
      ("01", "0110100100110101", "1111001000001100", "0111011100101001"), -- i=2877
      ("10", "0110100100110101", "1111001000001100", "0110000000000100"), -- i=2878
      ("11", "0110100100110101", "1111001000001100", "1111101100111101"), -- i=2879
      ("00", "0000111010100110", "1101101011011101", "1110100110000011"), -- i=2880
      ("01", "0000111010100110", "1101101011011101", "0011001111001001"), -- i=2881
      ("10", "0000111010100110", "1101101011011101", "0000101010000100"), -- i=2882
      ("11", "0000111010100110", "1101101011011101", "1101111011111111"), -- i=2883
      ("00", "1110111001111101", "0101100100110010", "0100011110101111"), -- i=2884
      ("01", "1110111001111101", "0101100100110010", "1001010101001011"), -- i=2885
      ("10", "1110111001111101", "0101100100110010", "0100100000110000"), -- i=2886
      ("11", "1110111001111101", "0101100100110010", "1111111101111111"), -- i=2887
      ("00", "0000000000001100", "1111011001100011", "1111011001101111"), -- i=2888
      ("01", "0000000000001100", "1111011001100011", "0000100110101001"), -- i=2889
      ("10", "0000000000001100", "1111011001100011", "0000000000000000"), -- i=2890
      ("11", "0000000000001100", "1111011001100011", "1111011001101111"), -- i=2891
      ("00", "1101001100011000", "1011101110001011", "1000111010100011"), -- i=2892
      ("01", "1101001100011000", "1011101110001011", "0001011110001101"), -- i=2893
      ("10", "1101001100011000", "1011101110001011", "1001001100001000"), -- i=2894
      ("11", "1101001100011000", "1011101110001011", "1111101110011011"), -- i=2895
      ("00", "1011110000010111", "0111110000010011", "0011100000101010"), -- i=2896
      ("01", "1011110000010111", "0111110000010011", "0100000000000100"), -- i=2897
      ("10", "1011110000010111", "0111110000010011", "0011110000010011"), -- i=2898
      ("11", "1011110000010111", "0111110000010011", "1111110000010111"), -- i=2899
      ("00", "1100100001111101", "0101101100000010", "0010001101111111"), -- i=2900
      ("01", "1100100001111101", "0101101100000010", "0110110101111011"), -- i=2901
      ("10", "1100100001111101", "0101101100000010", "0100100000000000"), -- i=2902
      ("11", "1100100001111101", "0101101100000010", "1101101101111111"), -- i=2903
      ("00", "1101101111001000", "0010100101100110", "0000010100101110"), -- i=2904
      ("01", "1101101111001000", "0010100101100110", "1011001001100010"), -- i=2905
      ("10", "1101101111001000", "0010100101100110", "0000100101000000"), -- i=2906
      ("11", "1101101111001000", "0010100101100110", "1111101111101110"), -- i=2907
      ("00", "0101100111101111", "0100000001100111", "1001101001010110"), -- i=2908
      ("01", "0101100111101111", "0100000001100111", "0001100110001000"), -- i=2909
      ("10", "0101100111101111", "0100000001100111", "0100000001100111"), -- i=2910
      ("11", "0101100111101111", "0100000001100111", "0101100111101111"), -- i=2911
      ("00", "0111011101000100", "1010111101011001", "0010011010011101"), -- i=2912
      ("01", "0111011101000100", "1010111101011001", "1100011111101011"), -- i=2913
      ("10", "0111011101000100", "1010111101011001", "0010011101000000"), -- i=2914
      ("11", "0111011101000100", "1010111101011001", "1111111101011101"), -- i=2915
      ("00", "1100100111000111", "0010000010100001", "1110101001101000"), -- i=2916
      ("01", "1100100111000111", "0010000010100001", "1010100100100110"), -- i=2917
      ("10", "1100100111000111", "0010000010100001", "0000000010000001"), -- i=2918
      ("11", "1100100111000111", "0010000010100001", "1110100111100111"), -- i=2919
      ("00", "0000000110110000", "1100111010001111", "1101000000111111"), -- i=2920
      ("01", "0000000110110000", "1100111010001111", "0011001100100001"), -- i=2921
      ("10", "0000000110110000", "1100111010001111", "0000000010000000"), -- i=2922
      ("11", "0000000110110000", "1100111010001111", "1100111110111111"), -- i=2923
      ("00", "1100011111000001", "1000111100000100", "0101011011000101"), -- i=2924
      ("01", "1100011111000001", "1000111100000100", "0011100010111101"), -- i=2925
      ("10", "1100011111000001", "1000111100000100", "1000011100000000"), -- i=2926
      ("11", "1100011111000001", "1000111100000100", "1100111111000101"), -- i=2927
      ("00", "0000010100111001", "0010000010111101", "0010010111110110"), -- i=2928
      ("01", "0000010100111001", "0010000010111101", "1110010001111100"), -- i=2929
      ("10", "0000010100111001", "0010000010111101", "0000000000111001"), -- i=2930
      ("11", "0000010100111001", "0010000010111101", "0010010110111101"), -- i=2931
      ("00", "0011101111100101", "1111001011100011", "0010111011001000"), -- i=2932
      ("01", "0011101111100101", "1111001011100011", "0100100100000010"), -- i=2933
      ("10", "0011101111100101", "1111001011100011", "0011001011100001"), -- i=2934
      ("11", "0011101111100101", "1111001011100011", "1111101111100111"), -- i=2935
      ("00", "1101101001111010", "1111111000101110", "1101100010101000"), -- i=2936
      ("01", "1101101001111010", "1111111000101110", "1101110001001100"), -- i=2937
      ("10", "1101101001111010", "1111111000101110", "1101101000101010"), -- i=2938
      ("11", "1101101001111010", "1111111000101110", "1111111001111110"), -- i=2939
      ("00", "0111101011110100", "1001000111101000", "0000110011011100"), -- i=2940
      ("01", "0111101011110100", "1001000111101000", "1110100100001100"), -- i=2941
      ("10", "0111101011110100", "1001000111101000", "0001000011100000"), -- i=2942
      ("11", "0111101011110100", "1001000111101000", "1111101111111100"), -- i=2943
      ("00", "1110001111001110", "0011110101100110", "0010000100110100"), -- i=2944
      ("01", "1110001111001110", "0011110101100110", "1010011001101000"), -- i=2945
      ("10", "1110001111001110", "0011110101100110", "0010000101000110"), -- i=2946
      ("11", "1110001111001110", "0011110101100110", "1111111111101110"), -- i=2947
      ("00", "0011101001100100", "0000001110110111", "0011111000011011"), -- i=2948
      ("01", "0011101001100100", "0000001110110111", "0011011010101101"), -- i=2949
      ("10", "0011101001100100", "0000001110110111", "0000001000100100"), -- i=2950
      ("11", "0011101001100100", "0000001110110111", "0011101111110111"), -- i=2951
      ("00", "1010101000110111", "1000001000110010", "0010110001101001"), -- i=2952
      ("01", "1010101000110111", "1000001000110010", "0010100000000101"), -- i=2953
      ("10", "1010101000110111", "1000001000110010", "1000001000110010"), -- i=2954
      ("11", "1010101000110111", "1000001000110010", "1010101000110111"), -- i=2955
      ("00", "1000001101010011", "1000111011101011", "0001001000111110"), -- i=2956
      ("01", "1000001101010011", "1000111011101011", "1111010001101000"), -- i=2957
      ("10", "1000001101010011", "1000111011101011", "1000001001000011"), -- i=2958
      ("11", "1000001101010011", "1000111011101011", "1000111111111011"), -- i=2959
      ("00", "0111011011010101", "0111000010101010", "1110011101111111"), -- i=2960
      ("01", "0111011011010101", "0111000010101010", "0000011000101011"), -- i=2961
      ("10", "0111011011010101", "0111000010101010", "0111000010000000"), -- i=2962
      ("11", "0111011011010101", "0111000010101010", "0111011011111111"), -- i=2963
      ("00", "1011010011110110", "0100001001110011", "1111011101101001"), -- i=2964
      ("01", "1011010011110110", "0100001001110011", "0111001010000011"), -- i=2965
      ("10", "1011010011110110", "0100001001110011", "0000000001110010"), -- i=2966
      ("11", "1011010011110110", "0100001001110011", "1111011011110111"), -- i=2967
      ("00", "1010100100110010", "0101111111110110", "0000100100101000"), -- i=2968
      ("01", "1010100100110010", "0101111111110110", "0100100100111100"), -- i=2969
      ("10", "1010100100110010", "0101111111110110", "0000100100110010"), -- i=2970
      ("11", "1010100100110010", "0101111111110110", "1111111111110110"), -- i=2971
      ("00", "0110000001111001", "0001100111011101", "0111101001010110"), -- i=2972
      ("01", "0110000001111001", "0001100111011101", "0100011010011100"), -- i=2973
      ("10", "0110000001111001", "0001100111011101", "0000000001011001"), -- i=2974
      ("11", "0110000001111001", "0001100111011101", "0111100111111101"), -- i=2975
      ("00", "0001011111010101", "0001011111011010", "0010111110101111"), -- i=2976
      ("01", "0001011111010101", "0001011111011010", "1111111111111011"), -- i=2977
      ("10", "0001011111010101", "0001011111011010", "0001011111010000"), -- i=2978
      ("11", "0001011111010101", "0001011111011010", "0001011111011111"), -- i=2979
      ("00", "0110100101010101", "0001111000010111", "1000011101101100"), -- i=2980
      ("01", "0110100101010101", "0001111000010111", "0100101100111110"), -- i=2981
      ("10", "0110100101010101", "0001111000010111", "0000100000010101"), -- i=2982
      ("11", "0110100101010101", "0001111000010111", "0111111101010111"), -- i=2983
      ("00", "0011110111010100", "1011101101001110", "1111100100100010"), -- i=2984
      ("01", "0011110111010100", "1011101101001110", "1000001010000110"), -- i=2985
      ("10", "0011110111010100", "1011101101001110", "0011100101000100"), -- i=2986
      ("11", "0011110111010100", "1011101101001110", "1011111111011110"), -- i=2987
      ("00", "0101111010000010", "0011111110100111", "1001111000101001"), -- i=2988
      ("01", "0101111010000010", "0011111110100111", "0001111011011011"), -- i=2989
      ("10", "0101111010000010", "0011111110100111", "0001111010000010"), -- i=2990
      ("11", "0101111010000010", "0011111110100111", "0111111110100111"), -- i=2991
      ("00", "1101010101100100", "0100000111000011", "0001011100100111"), -- i=2992
      ("01", "1101010101100100", "0100000111000011", "1001001110100001"), -- i=2993
      ("10", "1101010101100100", "0100000111000011", "0100000101000000"), -- i=2994
      ("11", "1101010101100100", "0100000111000011", "1101010111100111"), -- i=2995
      ("00", "0111001000001111", "1001101001111111", "0000110010001110"), -- i=2996
      ("01", "0111001000001111", "1001101001111111", "1101011110010000"), -- i=2997
      ("10", "0111001000001111", "1001101001111111", "0001001000001111"), -- i=2998
      ("11", "0111001000001111", "1001101001111111", "1111101001111111"), -- i=2999
      ("00", "1100010010100011", "1100011110111100", "1000110001011111"), -- i=3000
      ("01", "1100010010100011", "1100011110111100", "1111110011100111"), -- i=3001
      ("10", "1100010010100011", "1100011110111100", "1100010010100000"), -- i=3002
      ("11", "1100010010100011", "1100011110111100", "1100011110111111"), -- i=3003
      ("00", "1100111000011000", "1110111011010010", "1011110011101010"), -- i=3004
      ("01", "1100111000011000", "1110111011010010", "1101111101000110"), -- i=3005
      ("10", "1100111000011000", "1110111011010010", "1100111000010000"), -- i=3006
      ("11", "1100111000011000", "1110111011010010", "1110111011011010"), -- i=3007
      ("00", "1110111100001010", "1000111011100100", "0111110111101110"), -- i=3008
      ("01", "1110111100001010", "1000111011100100", "0110000000100110"), -- i=3009
      ("10", "1110111100001010", "1000111011100100", "1000111000000000"), -- i=3010
      ("11", "1110111100001010", "1000111011100100", "1110111111101110"), -- i=3011
      ("00", "0100011100010000", "0101110110010011", "1010010010100011"), -- i=3012
      ("01", "0100011100010000", "0101110110010011", "1110100101111101"), -- i=3013
      ("10", "0100011100010000", "0101110110010011", "0100010100010000"), -- i=3014
      ("11", "0100011100010000", "0101110110010011", "0101111110010011"), -- i=3015
      ("00", "1001001101010100", "1011110011011111", "0101000000110011"), -- i=3016
      ("01", "1001001101010100", "1011110011011111", "1101011001110101"), -- i=3017
      ("10", "1001001101010100", "1011110011011111", "1001000001010100"), -- i=3018
      ("11", "1001001101010100", "1011110011011111", "1011111111011111"), -- i=3019
      ("00", "1001010011010100", "1110001010010010", "0111011101100110"), -- i=3020
      ("01", "1001010011010100", "1110001010010010", "1011001001000010"), -- i=3021
      ("10", "1001010011010100", "1110001010010010", "1000000010010000"), -- i=3022
      ("11", "1001010011010100", "1110001010010010", "1111011011010110"), -- i=3023
      ("00", "0101101010111111", "1100011101010100", "0010001000010011"), -- i=3024
      ("01", "0101101010111111", "1100011101010100", "1001001101101011"), -- i=3025
      ("10", "0101101010111111", "1100011101010100", "0100001000010100"), -- i=3026
      ("11", "0101101010111111", "1100011101010100", "1101111111111111"), -- i=3027
      ("00", "0100110100010010", "1001100101011010", "1110011001101100"), -- i=3028
      ("01", "0100110100010010", "1001100101011010", "1011001110111000"), -- i=3029
      ("10", "0100110100010010", "1001100101011010", "0000100100010010"), -- i=3030
      ("11", "0100110100010010", "1001100101011010", "1101110101011010"), -- i=3031
      ("00", "0010001111110010", "0000001100011000", "0010011100001010"), -- i=3032
      ("01", "0010001111110010", "0000001100011000", "0010000011011010"), -- i=3033
      ("10", "0010001111110010", "0000001100011000", "0000001100010000"), -- i=3034
      ("11", "0010001111110010", "0000001100011000", "0010001111111010"), -- i=3035
      ("00", "1101001011101011", "1001010100111000", "0110100000100011"), -- i=3036
      ("01", "1101001011101011", "1001010100111000", "0011110110110011"), -- i=3037
      ("10", "1101001011101011", "1001010100111000", "1001000000101000"), -- i=3038
      ("11", "1101001011101011", "1001010100111000", "1101011111111011"), -- i=3039
      ("00", "1110000011111011", "1111101101011110", "1101110001011001"), -- i=3040
      ("01", "1110000011111011", "1111101101011110", "1110010110011101"), -- i=3041
      ("10", "1110000011111011", "1111101101011110", "1110000001011010"), -- i=3042
      ("11", "1110000011111011", "1111101101011110", "1111101111111111"), -- i=3043
      ("00", "0101000011010111", "1111100000010111", "0100100011101110"), -- i=3044
      ("01", "0101000011010111", "1111100000010111", "0101100011000000"), -- i=3045
      ("10", "0101000011010111", "1111100000010111", "0101000000010111"), -- i=3046
      ("11", "0101000011010111", "1111100000010111", "1111100011010111"), -- i=3047
      ("00", "1001010100010111", "0000110101011110", "1010001001110101"), -- i=3048
      ("01", "1001010100010111", "0000110101011110", "1000011110111001"), -- i=3049
      ("10", "1001010100010111", "0000110101011110", "0000010100010110"), -- i=3050
      ("11", "1001010100010111", "0000110101011110", "1001110101011111"), -- i=3051
      ("00", "1001101100111100", "1111111100100001", "1001101001011101"), -- i=3052
      ("01", "1001101100111100", "1111111100100001", "1001110000011011"), -- i=3053
      ("10", "1001101100111100", "1111111100100001", "1001101100100000"), -- i=3054
      ("11", "1001101100111100", "1111111100100001", "1111111100111101"), -- i=3055
      ("00", "1001110001010111", "0100001111010100", "1110000000101011"), -- i=3056
      ("01", "1001110001010111", "0100001111010100", "0101100010000011"), -- i=3057
      ("10", "1001110001010111", "0100001111010100", "0000000001010100"), -- i=3058
      ("11", "1001110001010111", "0100001111010100", "1101111111010111"), -- i=3059
      ("00", "1000101100111011", "1110111101000101", "0111101010000000"), -- i=3060
      ("01", "1000101100111011", "1110111101000101", "1001101111110110"), -- i=3061
      ("10", "1000101100111011", "1110111101000101", "1000101100000001"), -- i=3062
      ("11", "1000101100111011", "1110111101000101", "1110111101111111"), -- i=3063
      ("00", "1110110000111000", "1001010101001001", "1000000110000001"), -- i=3064
      ("01", "1110110000111000", "1001010101001001", "0101011011101111"), -- i=3065
      ("10", "1110110000111000", "1001010101001001", "1000010000001000"), -- i=3066
      ("11", "1110110000111000", "1001010101001001", "1111110101111001"), -- i=3067
      ("00", "1111101010100100", "0010011100010011", "0010000110110111"), -- i=3068
      ("01", "1111101010100100", "0010011100010011", "1101001110010001"), -- i=3069
      ("10", "1111101010100100", "0010011100010011", "0010001000000000"), -- i=3070
      ("11", "1111101010100100", "0010011100010011", "1111111110110111"), -- i=3071
      ("00", "1110100111001010", "0111011100010000", "0110000011011010"), -- i=3072
      ("01", "1110100111001010", "0111011100010000", "0111001010111010"), -- i=3073
      ("10", "1110100111001010", "0111011100010000", "0110000100000000"), -- i=3074
      ("11", "1110100111001010", "0111011100010000", "1111111111011010"), -- i=3075
      ("00", "0000101100010110", "0001111010010101", "0010100110101011"), -- i=3076
      ("01", "0000101100010110", "0001111010010101", "1110110010000001"), -- i=3077
      ("10", "0000101100010110", "0001111010010101", "0000101000010100"), -- i=3078
      ("11", "0000101100010110", "0001111010010101", "0001111110010111"), -- i=3079
      ("00", "1100011100001010", "0010111001010001", "1111010101011011"), -- i=3080
      ("01", "1100011100001010", "0010111001010001", "1001100010111001"), -- i=3081
      ("10", "1100011100001010", "0010111001010001", "0000011000000000"), -- i=3082
      ("11", "1100011100001010", "0010111001010001", "1110111101011011"), -- i=3083
      ("00", "1100101110110010", "1100100100010001", "1001010011000011"), -- i=3084
      ("01", "1100101110110010", "1100100100010001", "0000001010100001"), -- i=3085
      ("10", "1100101110110010", "1100100100010001", "1100100100010000"), -- i=3086
      ("11", "1100101110110010", "1100100100010001", "1100101110110011"), -- i=3087
      ("00", "0001011001110001", "0110011110101110", "0111111000011111"), -- i=3088
      ("01", "0001011001110001", "0110011110101110", "1010111011000011"), -- i=3089
      ("10", "0001011001110001", "0110011110101110", "0000011000100000"), -- i=3090
      ("11", "0001011001110001", "0110011110101110", "0111011111111111"), -- i=3091
      ("00", "1010000111111001", "1001111111011010", "0100000111010011"), -- i=3092
      ("01", "1010000111111001", "1001111111011010", "0000001000011111"), -- i=3093
      ("10", "1010000111111001", "1001111111011010", "1000000111011000"), -- i=3094
      ("11", "1010000111111001", "1001111111011010", "1011111111111011"), -- i=3095
      ("00", "0110100011110101", "0110010100111111", "1100111000110100"), -- i=3096
      ("01", "0110100011110101", "0110010100111111", "0000001110110110"), -- i=3097
      ("10", "0110100011110101", "0110010100111111", "0110000000110101"), -- i=3098
      ("11", "0110100011110101", "0110010100111111", "0110110111111111"), -- i=3099
      ("00", "0001001110101000", "1001100010100001", "1010110001001001"), -- i=3100
      ("01", "0001001110101000", "1001100010100001", "0111101100000111"), -- i=3101
      ("10", "0001001110101000", "1001100010100001", "0001000010100000"), -- i=3102
      ("11", "0001001110101000", "1001100010100001", "1001101110101001"), -- i=3103
      ("00", "0101011111101110", "1000000111111011", "1101100111101001"), -- i=3104
      ("01", "0101011111101110", "1000000111111011", "1101010111110011"), -- i=3105
      ("10", "0101011111101110", "1000000111111011", "0000000111101010"), -- i=3106
      ("11", "0101011111101110", "1000000111111011", "1101011111111111"), -- i=3107
      ("00", "1011000010111000", "0110110011101010", "0001110110100010"), -- i=3108
      ("01", "1011000010111000", "0110110011101010", "0100001111001110"), -- i=3109
      ("10", "1011000010111000", "0110110011101010", "0010000010101000"), -- i=3110
      ("11", "1011000010111000", "0110110011101010", "1111110011111010"), -- i=3111
      ("00", "0101000110100000", "1110000011010100", "0011001001110100"), -- i=3112
      ("01", "0101000110100000", "1110000011010100", "0111000011001100"), -- i=3113
      ("10", "0101000110100000", "1110000011010100", "0100000010000000"), -- i=3114
      ("11", "0101000110100000", "1110000011010100", "1111000111110100"), -- i=3115
      ("00", "1110010111010000", "1110001110001100", "1100100101011100"), -- i=3116
      ("01", "1110010111010000", "1110001110001100", "0000001001000100"), -- i=3117
      ("10", "1110010111010000", "1110001110001100", "1110000110000000"), -- i=3118
      ("11", "1110010111010000", "1110001110001100", "1110011111011100"), -- i=3119
      ("00", "1101110001011111", "1101110100001111", "1011100101101110"), -- i=3120
      ("01", "1101110001011111", "1101110100001111", "1111111101010000"), -- i=3121
      ("10", "1101110001011111", "1101110100001111", "1101110000001111"), -- i=3122
      ("11", "1101110001011111", "1101110100001111", "1101110101011111"), -- i=3123
      ("00", "0111000011001011", "0100000001110101", "1011000101000000"), -- i=3124
      ("01", "0111000011001011", "0100000001110101", "0011000001010110"), -- i=3125
      ("10", "0111000011001011", "0100000001110101", "0100000001000001"), -- i=3126
      ("11", "0111000011001011", "0100000001110101", "0111000011111111"), -- i=3127
      ("00", "1100100110001101", "0011100010100011", "0000001000110000"), -- i=3128
      ("01", "1100100110001101", "0011100010100011", "1001000011101010"), -- i=3129
      ("10", "1100100110001101", "0011100010100011", "0000100010000001"), -- i=3130
      ("11", "1100100110001101", "0011100010100011", "1111100110101111"), -- i=3131
      ("00", "0000101000101010", "1001101000000111", "1010010000110001"), -- i=3132
      ("01", "0000101000101010", "1001101000000111", "0111000000100011"), -- i=3133
      ("10", "0000101000101010", "1001101000000111", "0000101000000010"), -- i=3134
      ("11", "0000101000101010", "1001101000000111", "1001101000101111"), -- i=3135
      ("00", "1111111011100100", "0001010010100111", "0001001110001011"), -- i=3136
      ("01", "1111111011100100", "0001010010100111", "1110101000111101"), -- i=3137
      ("10", "1111111011100100", "0001010010100111", "0001010010100100"), -- i=3138
      ("11", "1111111011100100", "0001010010100111", "1111111011100111"), -- i=3139
      ("00", "1001011110000101", "1001011011001011", "0010111001010000"), -- i=3140
      ("01", "1001011110000101", "1001011011001011", "0000000010111010"), -- i=3141
      ("10", "1001011110000101", "1001011011001011", "1001011010000001"), -- i=3142
      ("11", "1001011110000101", "1001011011001011", "1001011111001111"), -- i=3143
      ("00", "0001000111001101", "0111011100100000", "1000100011101101"), -- i=3144
      ("01", "0001000111001101", "0111011100100000", "1001101010101101"), -- i=3145
      ("10", "0001000111001101", "0111011100100000", "0001000100000000"), -- i=3146
      ("11", "0001000111001101", "0111011100100000", "0111011111101101"), -- i=3147
      ("00", "1110010001100111", "0000000101011001", "1110010111000000"), -- i=3148
      ("01", "1110010001100111", "0000000101011001", "1110001100001110"), -- i=3149
      ("10", "1110010001100111", "0000000101011001", "0000000001000001"), -- i=3150
      ("11", "1110010001100111", "0000000101011001", "1110010101111111"), -- i=3151
      ("00", "1110110110111011", "1000000010101011", "0110111001100110"), -- i=3152
      ("01", "1110110110111011", "1000000010101011", "0110110100010000"), -- i=3153
      ("10", "1110110110111011", "1000000010101011", "1000000010101011"), -- i=3154
      ("11", "1110110110111011", "1000000010101011", "1110110110111011"), -- i=3155
      ("00", "0111000000011001", "1011001110011111", "0010001110111000"), -- i=3156
      ("01", "0111000000011001", "1011001110011111", "1011110001111010"), -- i=3157
      ("10", "0111000000011001", "1011001110011111", "0011000000011001"), -- i=3158
      ("11", "0111000000011001", "1011001110011111", "1111001110011111"), -- i=3159
      ("00", "0010001111000011", "0111101111100010", "1001111110100101"), -- i=3160
      ("01", "0010001111000011", "0111101111100010", "1010011111100001"), -- i=3161
      ("10", "0010001111000011", "0111101111100010", "0010001111000010"), -- i=3162
      ("11", "0010001111000011", "0111101111100010", "0111101111100011"), -- i=3163
      ("00", "0101100001000010", "1001010111110110", "1110111000111000"), -- i=3164
      ("01", "0101100001000010", "1001010111110110", "1100001001001100"), -- i=3165
      ("10", "0101100001000010", "1001010111110110", "0001000001000010"), -- i=3166
      ("11", "0101100001000010", "1001010111110110", "1101110111110110"), -- i=3167
      ("00", "0100111011110000", "1001111101101011", "1110111001011011"), -- i=3168
      ("01", "0100111011110000", "1001111101101011", "1010111110000101"), -- i=3169
      ("10", "0100111011110000", "1001111101101011", "0000111001100000"), -- i=3170
      ("11", "0100111011110000", "1001111101101011", "1101111111111011"), -- i=3171
      ("00", "1100100101111011", "1101000110110001", "1001101100101100"), -- i=3172
      ("01", "1100100101111011", "1101000110110001", "1111011111001010"), -- i=3173
      ("10", "1100100101111011", "1101000110110001", "1100000100110001"), -- i=3174
      ("11", "1100100101111011", "1101000110110001", "1101100111111011"), -- i=3175
      ("00", "0010111000000001", "1011001100011000", "1110000100011001"), -- i=3176
      ("01", "0010111000000001", "1011001100011000", "0111101011101001"), -- i=3177
      ("10", "0010111000000001", "1011001100011000", "0010001000000000"), -- i=3178
      ("11", "0010111000000001", "1011001100011000", "1011111100011001"), -- i=3179
      ("00", "1010100000100000", "1110001000000011", "1000101000100011"), -- i=3180
      ("01", "1010100000100000", "1110001000000011", "1100011000011101"), -- i=3181
      ("10", "1010100000100000", "1110001000000011", "1010000000000000"), -- i=3182
      ("11", "1010100000100000", "1110001000000011", "1110101000100011"), -- i=3183
      ("00", "1011000010100000", "1100011110001100", "0111100000101100"), -- i=3184
      ("01", "1011000010100000", "1100011110001100", "1110100100010100"), -- i=3185
      ("10", "1011000010100000", "1100011110001100", "1000000010000000"), -- i=3186
      ("11", "1011000010100000", "1100011110001100", "1111011110101100"), -- i=3187
      ("00", "0101010100001100", "1110000101111001", "0011011010000101"), -- i=3188
      ("01", "0101010100001100", "1110000101111001", "0111001110010011"), -- i=3189
      ("10", "0101010100001100", "1110000101111001", "0100000100001000"), -- i=3190
      ("11", "0101010100001100", "1110000101111001", "1111010101111101"), -- i=3191
      ("00", "0011101100110010", "1101011100110110", "0001001001101000"), -- i=3192
      ("01", "0011101100110010", "1101011100110110", "0110001111111100"), -- i=3193
      ("10", "0011101100110010", "1101011100110110", "0001001100110010"), -- i=3194
      ("11", "0011101100110010", "1101011100110110", "1111111100110110"), -- i=3195
      ("00", "1000101100001101", "0100110101011100", "1101100001101001"), -- i=3196
      ("01", "1000101100001101", "0100110101011100", "0011110110110001"), -- i=3197
      ("10", "1000101100001101", "0100110101011100", "0000100100001100"), -- i=3198
      ("11", "1000101100001101", "0100110101011100", "1100111101011101"), -- i=3199
      ("00", "1101000111010010", "0111011010110011", "0100100010000101"), -- i=3200
      ("01", "1101000111010010", "0111011010110011", "0101101100011111"), -- i=3201
      ("10", "1101000111010010", "0111011010110011", "0101000010010010"), -- i=3202
      ("11", "1101000111010010", "0111011010110011", "1111011111110011"), -- i=3203
      ("00", "0101001100100110", "0111101110111110", "1100111011100100"), -- i=3204
      ("01", "0101001100100110", "0111101110111110", "1101011101101000"), -- i=3205
      ("10", "0101001100100110", "0111101110111110", "0101001100100110"), -- i=3206
      ("11", "0101001100100110", "0111101110111110", "0111101110111110"), -- i=3207
      ("00", "1011000000011111", "1011000111010010", "0110000111110001"), -- i=3208
      ("01", "1011000000011111", "1011000111010010", "1111111001001101"), -- i=3209
      ("10", "1011000000011111", "1011000111010010", "1011000000010010"), -- i=3210
      ("11", "1011000000011111", "1011000111010010", "1011000111011111"), -- i=3211
      ("00", "1111011100001110", "0010110000000010", "0010001100010000"), -- i=3212
      ("01", "1111011100001110", "0010110000000010", "1100101100001100"), -- i=3213
      ("10", "1111011100001110", "0010110000000010", "0010010000000010"), -- i=3214
      ("11", "1111011100001110", "0010110000000010", "1111111100001110"), -- i=3215
      ("00", "0001000011100011", "1101000111010111", "1110001010111010"), -- i=3216
      ("01", "0001000011100011", "1101000111010111", "0011111100001100"), -- i=3217
      ("10", "0001000011100011", "1101000111010111", "0001000011000011"), -- i=3218
      ("11", "0001000011100011", "1101000111010111", "1101000111110111"), -- i=3219
      ("00", "1010101001101100", "1110110100100011", "1001011110001111"), -- i=3220
      ("01", "1010101001101100", "1110110100100011", "1011110101001001"), -- i=3221
      ("10", "1010101001101100", "1110110100100011", "1010100000100000"), -- i=3222
      ("11", "1010101001101100", "1110110100100011", "1110111101101111"), -- i=3223
      ("00", "1000110111000101", "0001000010110100", "1001111001111001"), -- i=3224
      ("01", "1000110111000101", "0001000010110100", "0111110100010001"), -- i=3225
      ("10", "1000110111000101", "0001000010110100", "0000000010000100"), -- i=3226
      ("11", "1000110111000101", "0001000010110100", "1001110111110101"), -- i=3227
      ("00", "0101110010111111", "1001000000001000", "1110110011000111"), -- i=3228
      ("01", "0101110010111111", "1001000000001000", "1100110010110111"), -- i=3229
      ("10", "0101110010111111", "1001000000001000", "0001000000001000"), -- i=3230
      ("11", "0101110010111111", "1001000000001000", "1101110010111111"), -- i=3231
      ("00", "1000110010000101", "0010110001010000", "1011100011010101"), -- i=3232
      ("01", "1000110010000101", "0010110001010000", "0110000000110101"), -- i=3233
      ("10", "1000110010000101", "0010110001010000", "0000110000000000"), -- i=3234
      ("11", "1000110010000101", "0010110001010000", "1010110011010101"), -- i=3235
      ("00", "1100011011111101", "0111111110101010", "0100011010100111"), -- i=3236
      ("01", "1100011011111101", "0111111110101010", "0100011101010011"), -- i=3237
      ("10", "1100011011111101", "0111111110101010", "0100011010101000"), -- i=3238
      ("11", "1100011011111101", "0111111110101010", "1111111111111111"), -- i=3239
      ("00", "1010010001111011", "0110010000100000", "0000100010011011"), -- i=3240
      ("01", "1010010001111011", "0110010000100000", "0100000001011011"), -- i=3241
      ("10", "1010010001111011", "0110010000100000", "0010010000100000"), -- i=3242
      ("11", "1010010001111011", "0110010000100000", "1110010001111011"), -- i=3243
      ("00", "0101000101001110", "1010001111100111", "1111010100110101"), -- i=3244
      ("01", "0101000101001110", "1010001111100111", "1010110101100111"), -- i=3245
      ("10", "0101000101001110", "1010001111100111", "0000000101000110"), -- i=3246
      ("11", "0101000101001110", "1010001111100111", "1111001111101111"), -- i=3247
      ("00", "1100010001010001", "1010101010011001", "0110111011101010"), -- i=3248
      ("01", "1100010001010001", "1010101010011001", "0001100110111000"), -- i=3249
      ("10", "1100010001010001", "1010101010011001", "1000000000010001"), -- i=3250
      ("11", "1100010001010001", "1010101010011001", "1110111011011001"), -- i=3251
      ("00", "1101111001110100", "0110011100101000", "0100010110011100"), -- i=3252
      ("01", "1101111001110100", "0110011100101000", "0111011101001100"), -- i=3253
      ("10", "1101111001110100", "0110011100101000", "0100011000100000"), -- i=3254
      ("11", "1101111001110100", "0110011100101000", "1111111101111100"), -- i=3255
      ("00", "0010010100110100", "1011101101001111", "1110000010000011"), -- i=3256
      ("01", "0010010100110100", "1011101101001111", "0110100111100101"), -- i=3257
      ("10", "0010010100110100", "1011101101001111", "0010000100000100"), -- i=3258
      ("11", "0010010100110100", "1011101101001111", "1011111101111111"), -- i=3259
      ("00", "1110001111000011", "1001001001010101", "0111011000011000"), -- i=3260
      ("01", "1110001111000011", "1001001001010101", "0101000101101110"), -- i=3261
      ("10", "1110001111000011", "1001001001010101", "1000001001000001"), -- i=3262
      ("11", "1110001111000011", "1001001001010101", "1111001111010111"), -- i=3263
      ("00", "1100010111110100", "0101010111000000", "0001101110110100"), -- i=3264
      ("01", "1100010111110100", "0101010111000000", "0111000000110100"), -- i=3265
      ("10", "1100010111110100", "0101010111000000", "0100010111000000"), -- i=3266
      ("11", "1100010111110100", "0101010111000000", "1101010111110100"), -- i=3267
      ("00", "0111010110111010", "1111010110101111", "0110101101101001"), -- i=3268
      ("01", "0111010110111010", "1111010110101111", "1000000000001011"), -- i=3269
      ("10", "0111010110111010", "1111010110101111", "0111010110101010"), -- i=3270
      ("11", "0111010110111010", "1111010110101111", "1111010110111111"), -- i=3271
      ("00", "0011110111001111", "0001010000011100", "0101000111101011"), -- i=3272
      ("01", "0011110111001111", "0001010000011100", "0010100110110011"), -- i=3273
      ("10", "0011110111001111", "0001010000011100", "0001010000001100"), -- i=3274
      ("11", "0011110111001111", "0001010000011100", "0011110111011111"), -- i=3275
      ("00", "0001101010100000", "0100000010000100", "0101101100100100"), -- i=3276
      ("01", "0001101010100000", "0100000010000100", "1101101000011100"), -- i=3277
      ("10", "0001101010100000", "0100000010000100", "0000000010000000"), -- i=3278
      ("11", "0001101010100000", "0100000010000100", "0101101010100100"), -- i=3279
      ("00", "0011001111100100", "0011010010010010", "0110100001110110"), -- i=3280
      ("01", "0011001111100100", "0011010010010010", "1111111101010010"), -- i=3281
      ("10", "0011001111100100", "0011010010010010", "0011000010000000"), -- i=3282
      ("11", "0011001111100100", "0011010010010010", "0011011111110110"), -- i=3283
      ("00", "0100010110110011", "1111110011101001", "0100001010011100"), -- i=3284
      ("01", "0100010110110011", "1111110011101001", "0100100011001010"), -- i=3285
      ("10", "0100010110110011", "1111110011101001", "0100010010100001"), -- i=3286
      ("11", "0100010110110011", "1111110011101001", "1111110111111011"), -- i=3287
      ("00", "1010110101111101", "0011001011101000", "1110000001100101"), -- i=3288
      ("01", "1010110101111101", "0011001011101000", "0111101010010101"), -- i=3289
      ("10", "1010110101111101", "0011001011101000", "0010000001101000"), -- i=3290
      ("11", "1010110101111101", "0011001011101000", "1011111111111101"), -- i=3291
      ("00", "0101011011010011", "0101111111011001", "1011011010101100"), -- i=3292
      ("01", "0101011011010011", "0101111111011001", "1111011011111010"), -- i=3293
      ("10", "0101011011010011", "0101111111011001", "0101011011010001"), -- i=3294
      ("11", "0101011011010011", "0101111111011001", "0101111111011011"), -- i=3295
      ("00", "1011001010110111", "0011111101110101", "1111001000101100"), -- i=3296
      ("01", "1011001010110111", "0011111101110101", "0111001101000010"), -- i=3297
      ("10", "1011001010110111", "0011111101110101", "0011001000110101"), -- i=3298
      ("11", "1011001010110111", "0011111101110101", "1011111111110111"), -- i=3299
      ("00", "1101101110110110", "1000000101101110", "0101110100100100"), -- i=3300
      ("01", "1101101110110110", "1000000101101110", "0101101001001000"), -- i=3301
      ("10", "1101101110110110", "1000000101101110", "1000000100100110"), -- i=3302
      ("11", "1101101110110110", "1000000101101110", "1101101111111110"), -- i=3303
      ("00", "0111111000111011", "0111011110110001", "1111010111101100"), -- i=3304
      ("01", "0111111000111011", "0111011110110001", "0000011010001010"), -- i=3305
      ("10", "0111111000111011", "0111011110110001", "0111011000110001"), -- i=3306
      ("11", "0111111000111011", "0111011110110001", "0111111110111011"), -- i=3307
      ("00", "1001100011111111", "1001110000011001", "0011010100011000"), -- i=3308
      ("01", "1001100011111111", "1001110000011001", "1111110011100110"), -- i=3309
      ("10", "1001100011111111", "1001110000011001", "1001100000011001"), -- i=3310
      ("11", "1001100011111111", "1001110000011001", "1001110011111111"), -- i=3311
      ("00", "1000101000000001", "0100001111111011", "1100110111111100"), -- i=3312
      ("01", "1000101000000001", "0100001111111011", "0100011000000110"), -- i=3313
      ("10", "1000101000000001", "0100001111111011", "0000001000000001"), -- i=3314
      ("11", "1000101000000001", "0100001111111011", "1100101111111011"), -- i=3315
      ("00", "1001001011100001", "0010010100000101", "1011011111100110"), -- i=3316
      ("01", "1001001011100001", "0010010100000101", "0110110111011100"), -- i=3317
      ("10", "1001001011100001", "0010010100000101", "0000000000000001"), -- i=3318
      ("11", "1001001011100001", "0010010100000101", "1011011111100101"), -- i=3319
      ("00", "0101000001011110", "0110010101010111", "1011010110110101"), -- i=3320
      ("01", "0101000001011110", "0110010101010111", "1110101100000111"), -- i=3321
      ("10", "0101000001011110", "0110010101010111", "0100000001010110"), -- i=3322
      ("11", "0101000001011110", "0110010101010111", "0111010101011111"), -- i=3323
      ("00", "1110011000010010", "1110101100001000", "1101000100011010"), -- i=3324
      ("01", "1110011000010010", "1110101100001000", "1111101100001010"), -- i=3325
      ("10", "1110011000010010", "1110101100001000", "1110001000000000"), -- i=3326
      ("11", "1110011000010010", "1110101100001000", "1110111100011010"), -- i=3327
      ("00", "1000010111001110", "0000110100100100", "1001001011110010"), -- i=3328
      ("01", "1000010111001110", "0000110100100100", "0111100010101010"), -- i=3329
      ("10", "1000010111001110", "0000110100100100", "0000010100000100"), -- i=3330
      ("11", "1000010111001110", "0000110100100100", "1000110111101110"), -- i=3331
      ("00", "1100001100111110", "1110110011011110", "1011000000011100"), -- i=3332
      ("01", "1100001100111110", "1110110011011110", "1101011001100000"), -- i=3333
      ("10", "1100001100111110", "1110110011011110", "1100000000011110"), -- i=3334
      ("11", "1100001100111110", "1110110011011110", "1110111111111110"), -- i=3335
      ("00", "1110010100111001", "1101000000100011", "1011010101011100"), -- i=3336
      ("01", "1110010100111001", "1101000000100011", "0001010100010110"), -- i=3337
      ("10", "1110010100111001", "1101000000100011", "1100000000100001"), -- i=3338
      ("11", "1110010100111001", "1101000000100011", "1111010100111011"), -- i=3339
      ("00", "0100100000111011", "0100001001111100", "1000101010110111"), -- i=3340
      ("01", "0100100000111011", "0100001001111100", "0000010110111111"), -- i=3341
      ("10", "0100100000111011", "0100001001111100", "0100000000111000"), -- i=3342
      ("11", "0100100000111011", "0100001001111100", "0100101001111111"), -- i=3343
      ("00", "0110010110101111", "0110010101010110", "1100101100000101"), -- i=3344
      ("01", "0110010110101111", "0110010101010110", "0000000001011001"), -- i=3345
      ("10", "0110010110101111", "0110010101010110", "0110010100000110"), -- i=3346
      ("11", "0110010110101111", "0110010101010110", "0110010111111111"), -- i=3347
      ("00", "0100001110111010", "0100100011000010", "1000110001111100"), -- i=3348
      ("01", "0100001110111010", "0100100011000010", "1111101011111000"), -- i=3349
      ("10", "0100001110111010", "0100100011000010", "0100000010000010"), -- i=3350
      ("11", "0100001110111010", "0100100011000010", "0100101111111010"), -- i=3351
      ("00", "1101010111001111", "1110100001110010", "1011111001000001"), -- i=3352
      ("01", "1101010111001111", "1110100001110010", "1110110101011101"), -- i=3353
      ("10", "1101010111001111", "1110100001110010", "1100000001000010"), -- i=3354
      ("11", "1101010111001111", "1110100001110010", "1111110111111111"), -- i=3355
      ("00", "0010100100100110", "0011100111100011", "0110001100001001"), -- i=3356
      ("01", "0010100100100110", "0011100111100011", "1110111101000011"), -- i=3357
      ("10", "0010100100100110", "0011100111100011", "0010100100100010"), -- i=3358
      ("11", "0010100100100110", "0011100111100011", "0011100111100111"), -- i=3359
      ("00", "0110011001011000", "1100011100001011", "0010110101100011"), -- i=3360
      ("01", "0110011001011000", "1100011100001011", "1001111101001101"), -- i=3361
      ("10", "0110011001011000", "1100011100001011", "0100011000001000"), -- i=3362
      ("11", "0110011001011000", "1100011100001011", "1110011101011011"), -- i=3363
      ("00", "1001101111110100", "1000000000110001", "0001110000100101"), -- i=3364
      ("01", "1001101111110100", "1000000000110001", "0001101111000011"), -- i=3365
      ("10", "1001101111110100", "1000000000110001", "1000000000110000"), -- i=3366
      ("11", "1001101111110100", "1000000000110001", "1001101111110101"), -- i=3367
      ("00", "1010001010011100", "1001011010011111", "0011100100111011"), -- i=3368
      ("01", "1010001010011100", "1001011010011111", "0000101111111101"), -- i=3369
      ("10", "1010001010011100", "1001011010011111", "1000001010011100"), -- i=3370
      ("11", "1010001010011100", "1001011010011111", "1011011010011111"), -- i=3371
      ("00", "0000001010010111", "0101110001000001", "0101111011011000"), -- i=3372
      ("01", "0000001010010111", "0101110001000001", "1010011001010110"), -- i=3373
      ("10", "0000001010010111", "0101110001000001", "0000000000000001"), -- i=3374
      ("11", "0000001010010111", "0101110001000001", "0101111011010111"), -- i=3375
      ("00", "1011001011010011", "1101000100110000", "1000010000000011"), -- i=3376
      ("01", "1011001011010011", "1101000100110000", "1110000110100011"), -- i=3377
      ("10", "1011001011010011", "1101000100110000", "1001000000010000"), -- i=3378
      ("11", "1011001011010011", "1101000100110000", "1111001111110011"), -- i=3379
      ("00", "1000001011011010", "1110101001111011", "0110110101010101"), -- i=3380
      ("01", "1000001011011010", "1110101001111011", "1001100001011111"), -- i=3381
      ("10", "1000001011011010", "1110101001111011", "1000001001011010"), -- i=3382
      ("11", "1000001011011010", "1110101001111011", "1110101011111011"), -- i=3383
      ("00", "1000100101111001", "1101110100011010", "0110011010010011"), -- i=3384
      ("01", "1000100101111001", "1101110100011010", "1010110001011111"), -- i=3385
      ("10", "1000100101111001", "1101110100011010", "1000100100011000"), -- i=3386
      ("11", "1000100101111001", "1101110100011010", "1101110101111011"), -- i=3387
      ("00", "1010001001010011", "0010111110011110", "1101000111110001"), -- i=3388
      ("01", "1010001001010011", "0010111110011110", "0111001010110101"), -- i=3389
      ("10", "1010001001010011", "0010111110011110", "0010001000010010"), -- i=3390
      ("11", "1010001001010011", "0010111110011110", "1010111111011111"), -- i=3391
      ("00", "1100101001001100", "1101010000111100", "1001111010001000"), -- i=3392
      ("01", "1100101001001100", "1101010000111100", "1111011000010000"), -- i=3393
      ("10", "1100101001001100", "1101010000111100", "1100000000001100"), -- i=3394
      ("11", "1100101001001100", "1101010000111100", "1101111001111100"), -- i=3395
      ("00", "1000011100100100", "1001011011000100", "0001110111101000"), -- i=3396
      ("01", "1000011100100100", "1001011011000100", "1111000001100000"), -- i=3397
      ("10", "1000011100100100", "1001011011000100", "1000011000000100"), -- i=3398
      ("11", "1000011100100100", "1001011011000100", "1001011111100100"), -- i=3399
      ("00", "1100111010000111", "0011010110111100", "0000010001000011"), -- i=3400
      ("01", "1100111010000111", "0011010110111100", "1001100011001011"), -- i=3401
      ("10", "1100111010000111", "0011010110111100", "0000010010000100"), -- i=3402
      ("11", "1100111010000111", "0011010110111100", "1111111110111111"), -- i=3403
      ("00", "0111111001011110", "0011011011101000", "1011010101000110"), -- i=3404
      ("01", "0111111001011110", "0011011011101000", "0100011101110110"), -- i=3405
      ("10", "0111111001011110", "0011011011101000", "0011011001001000"), -- i=3406
      ("11", "0111111001011110", "0011011011101000", "0111111011111110"), -- i=3407
      ("00", "0010011101101001", "0000110011110011", "0011010001011100"), -- i=3408
      ("01", "0010011101101001", "0000110011110011", "0001101001110110"), -- i=3409
      ("10", "0010011101101001", "0000110011110011", "0000010001100001"), -- i=3410
      ("11", "0010011101101001", "0000110011110011", "0010111111111011"), -- i=3411
      ("00", "1111111010010101", "0100100100000111", "0100011110011100"), -- i=3412
      ("01", "1111111010010101", "0100100100000111", "1011010110001110"), -- i=3413
      ("10", "1111111010010101", "0100100100000111", "0100100000000101"), -- i=3414
      ("11", "1111111010010101", "0100100100000111", "1111111110010111"), -- i=3415
      ("00", "0110010100111000", "0001111101000100", "1000010001111100"), -- i=3416
      ("01", "0110010100111000", "0001111101000100", "0100010111110100"), -- i=3417
      ("10", "0110010100111000", "0001111101000100", "0000010100000000"), -- i=3418
      ("11", "0110010100111000", "0001111101000100", "0111111101111100"), -- i=3419
      ("00", "1101011010010001", "0111001101001110", "0100100111011111"), -- i=3420
      ("01", "1101011010010001", "0111001101001110", "0110001101000011"), -- i=3421
      ("10", "1101011010010001", "0111001101001110", "0101001000000000"), -- i=3422
      ("11", "1101011010010001", "0111001101001110", "1111011111011111"), -- i=3423
      ("00", "1011011000111010", "0110000111101001", "0001100000100011"), -- i=3424
      ("01", "1011011000111010", "0110000111101001", "0101010001010001"), -- i=3425
      ("10", "1011011000111010", "0110000111101001", "0010000000101000"), -- i=3426
      ("11", "1011011000111010", "0110000111101001", "1111011111111011"), -- i=3427
      ("00", "1001100100100000", "1111000100000011", "1000101000100011"), -- i=3428
      ("01", "1001100100100000", "1111000100000011", "1010100000011101"), -- i=3429
      ("10", "1001100100100000", "1111000100000011", "1001000100000000"), -- i=3430
      ("11", "1001100100100000", "1111000100000011", "1111100100100011"), -- i=3431
      ("00", "0010011001100111", "0101000000001110", "0111011001110101"), -- i=3432
      ("01", "0010011001100111", "0101000000001110", "1101011001011001"), -- i=3433
      ("10", "0010011001100111", "0101000000001110", "0000000000000110"), -- i=3434
      ("11", "0010011001100111", "0101000000001110", "0111011001101111"), -- i=3435
      ("00", "1010000001111110", "0010101000000110", "1100101010000100"), -- i=3436
      ("01", "1010000001111110", "0010101000000110", "0111011001111000"), -- i=3437
      ("10", "1010000001111110", "0010101000000110", "0010000000000110"), -- i=3438
      ("11", "1010000001111110", "0010101000000110", "1010101001111110"), -- i=3439
      ("00", "1110010110111111", "1011100010101011", "1001111001101010"), -- i=3440
      ("01", "1110010110111111", "1011100010101011", "0010110100010100"), -- i=3441
      ("10", "1110010110111111", "1011100010101011", "1010000010101011"), -- i=3442
      ("11", "1110010110111111", "1011100010101011", "1111110110111111"), -- i=3443
      ("00", "0011010011010010", "0000000000100011", "0011010011110101"), -- i=3444
      ("01", "0011010011010010", "0000000000100011", "0011010010101111"), -- i=3445
      ("10", "0011010011010010", "0000000000100011", "0000000000000010"), -- i=3446
      ("11", "0011010011010010", "0000000000100011", "0011010011110011"), -- i=3447
      ("00", "0000000010001010", "0100001100000001", "0100001110001011"), -- i=3448
      ("01", "0000000010001010", "0100001100000001", "1011110110001001"), -- i=3449
      ("10", "0000000010001010", "0100001100000001", "0000000000000000"), -- i=3450
      ("11", "0000000010001010", "0100001100000001", "0100001110001011"), -- i=3451
      ("00", "0111101010101100", "1111001110010010", "0110111000111110"), -- i=3452
      ("01", "0111101010101100", "1111001110010010", "1000011100011010"), -- i=3453
      ("10", "0111101010101100", "1111001110010010", "0111001010000000"), -- i=3454
      ("11", "0111101010101100", "1111001110010010", "1111101110111110"), -- i=3455
      ("00", "0110000111111101", "0011011110101011", "1001100110101000"), -- i=3456
      ("01", "0110000111111101", "0011011110101011", "0010101001010010"), -- i=3457
      ("10", "0110000111111101", "0011011110101011", "0010000110101001"), -- i=3458
      ("11", "0110000111111101", "0011011110101011", "0111011111111111"), -- i=3459
      ("00", "1100111110011010", "0100001101010111", "0001001011110001"), -- i=3460
      ("01", "1100111110011010", "0100001101010111", "1000110001000011"), -- i=3461
      ("10", "1100111110011010", "0100001101010111", "0100001100010010"), -- i=3462
      ("11", "1100111110011010", "0100001101010111", "1100111111011111"), -- i=3463
      ("00", "1100111011101111", "0001001110101001", "1110001010011000"), -- i=3464
      ("01", "1100111011101111", "0001001110101001", "1011101101000110"), -- i=3465
      ("10", "1100111011101111", "0001001110101001", "0000001010101001"), -- i=3466
      ("11", "1100111011101111", "0001001110101001", "1101111111101111"), -- i=3467
      ("00", "0010010000100110", "0101100101101101", "0111110110010011"), -- i=3468
      ("01", "0010010000100110", "0101100101101101", "1100101010111001"), -- i=3469
      ("10", "0010010000100110", "0101100101101101", "0000000000100100"), -- i=3470
      ("11", "0010010000100110", "0101100101101101", "0111110101101111"), -- i=3471
      ("00", "1100001110101101", "0000100111010010", "1100110101111111"), -- i=3472
      ("01", "1100001110101101", "0000100111010010", "1011100111011011"), -- i=3473
      ("10", "1100001110101101", "0000100111010010", "0000000110000000"), -- i=3474
      ("11", "1100001110101101", "0000100111010010", "1100101111111111"), -- i=3475
      ("00", "1011001111100011", "0010010111011110", "1101100111000001"), -- i=3476
      ("01", "1011001111100011", "0010010111011110", "1000111000000101"), -- i=3477
      ("10", "1011001111100011", "0010010111011110", "0010000111000010"), -- i=3478
      ("11", "1011001111100011", "0010010111011110", "1011011111111111"), -- i=3479
      ("00", "1100010100010100", "1101111010001101", "1010001110100001"), -- i=3480
      ("01", "1100010100010100", "1101111010001101", "1110011010000111"), -- i=3481
      ("10", "1100010100010100", "1101111010001101", "1100010000000100"), -- i=3482
      ("11", "1100010100010100", "1101111010001101", "1101111110011101"), -- i=3483
      ("00", "0011010101011100", "1000011100111001", "1011110010010101"), -- i=3484
      ("01", "0011010101011100", "1000011100111001", "1010111000100011"), -- i=3485
      ("10", "0011010101011100", "1000011100111001", "0000010100011000"), -- i=3486
      ("11", "0011010101011100", "1000011100111001", "1011011101111101"), -- i=3487
      ("00", "1100001001111010", "0111100011001111", "0011101101001001"), -- i=3488
      ("01", "1100001001111010", "0111100011001111", "0100100110101011"), -- i=3489
      ("10", "1100001001111010", "0111100011001111", "0100000001001010"), -- i=3490
      ("11", "1100001001111010", "0111100011001111", "1111101011111111"), -- i=3491
      ("00", "0011110011111101", "1000001000001101", "1011111100001010"), -- i=3492
      ("01", "0011110011111101", "1000001000001101", "1011101011110000"), -- i=3493
      ("10", "0011110011111101", "1000001000001101", "0000000000001101"), -- i=3494
      ("11", "0011110011111101", "1000001000001101", "1011111011111101"), -- i=3495
      ("00", "1001101100010001", "0001101010110001", "1011010111000010"), -- i=3496
      ("01", "1001101100010001", "0001101010110001", "1000000001100000"), -- i=3497
      ("10", "1001101100010001", "0001101010110001", "0001101000010001"), -- i=3498
      ("11", "1001101100010001", "0001101010110001", "1001101110110001"), -- i=3499
      ("00", "0001011101011011", "1101010001010110", "1110101110110001"), -- i=3500
      ("01", "0001011101011011", "1101010001010110", "0100001100000101"), -- i=3501
      ("10", "0001011101011011", "1101010001010110", "0001010001010010"), -- i=3502
      ("11", "0001011101011011", "1101010001010110", "1101011101011111"), -- i=3503
      ("00", "1011011011010010", "0111001100011001", "0010100111101011"), -- i=3504
      ("01", "1011011011010010", "0111001100011001", "0100001110111001"), -- i=3505
      ("10", "1011011011010010", "0111001100011001", "0011001000010000"), -- i=3506
      ("11", "1011011011010010", "0111001100011001", "1111011111011011"), -- i=3507
      ("00", "1101000001100010", "0110010100000001", "0011010101100011"), -- i=3508
      ("01", "1101000001100010", "0110010100000001", "0110101101100001"), -- i=3509
      ("10", "1101000001100010", "0110010100000001", "0100000000000000"), -- i=3510
      ("11", "1101000001100010", "0110010100000001", "1111010101100011"), -- i=3511
      ("00", "1110100000010100", "1010000101010100", "1000100101101000"), -- i=3512
      ("01", "1110100000010100", "1010000101010100", "0100011011000000"), -- i=3513
      ("10", "1110100000010100", "1010000101010100", "1010000000010100"), -- i=3514
      ("11", "1110100000010100", "1010000101010100", "1110100101010100"), -- i=3515
      ("00", "0111011001011010", "0010101011110011", "1010000101001101"), -- i=3516
      ("01", "0111011001011010", "0010101011110011", "0100101101100111"), -- i=3517
      ("10", "0111011001011010", "0010101011110011", "0010001001010010"), -- i=3518
      ("11", "0111011001011010", "0010101011110011", "0111111011111011"), -- i=3519
      ("00", "0111100001010110", "1101001010011110", "0100101011110100"), -- i=3520
      ("01", "0111100001010110", "1101001010011110", "1010010110111000"), -- i=3521
      ("10", "0111100001010110", "1101001010011110", "0101000000010110"), -- i=3522
      ("11", "0111100001010110", "1101001010011110", "1111101011011110"), -- i=3523
      ("00", "1110100011001000", "0110101001000110", "0101001100001110"), -- i=3524
      ("01", "1110100011001000", "0110101001000110", "0111111010000010"), -- i=3525
      ("10", "1110100011001000", "0110101001000110", "0110100001000000"), -- i=3526
      ("11", "1110100011001000", "0110101001000110", "1110101011001110"), -- i=3527
      ("00", "0101011111110110", "0101100011011110", "1011000011010100"), -- i=3528
      ("01", "0101011111110110", "0101100011011110", "1111111100011000"), -- i=3529
      ("10", "0101011111110110", "0101100011011110", "0101000011010110"), -- i=3530
      ("11", "0101011111110110", "0101100011011110", "0101111111111110"), -- i=3531
      ("00", "1010110010010101", "1001000110010000", "0011111000100101"), -- i=3532
      ("01", "1010110010010101", "1001000110010000", "0001101100000101"), -- i=3533
      ("10", "1010110010010101", "1001000110010000", "1000000010010000"), -- i=3534
      ("11", "1010110010010101", "1001000110010000", "1011110110010101"), -- i=3535
      ("00", "1110010111001100", "1111100100110001", "1101111011111101"), -- i=3536
      ("01", "1110010111001100", "1111100100110001", "1110110010011011"), -- i=3537
      ("10", "1110010111001100", "1111100100110001", "1110000100000000"), -- i=3538
      ("11", "1110010111001100", "1111100100110001", "1111110111111101"), -- i=3539
      ("00", "0101000000001010", "1001010001111001", "1110010010000011"), -- i=3540
      ("01", "0101000000001010", "1001010001111001", "1011101110010001"), -- i=3541
      ("10", "0101000000001010", "1001010001111001", "0001000000001000"), -- i=3542
      ("11", "0101000000001010", "1001010001111001", "1101010001111011"), -- i=3543
      ("00", "1010100011011110", "1011011111111111", "0110000011011101"), -- i=3544
      ("01", "1010100011011110", "1011011111111111", "1111000011011111"), -- i=3545
      ("10", "1010100011011110", "1011011111111111", "1010000011011110"), -- i=3546
      ("11", "1010100011011110", "1011011111111111", "1011111111111111"), -- i=3547
      ("00", "1110001010000010", "0101101111110101", "0011111001110111"), -- i=3548
      ("01", "1110001010000010", "0101101111110101", "1000011010001101"), -- i=3549
      ("10", "1110001010000010", "0101101111110101", "0100001010000000"), -- i=3550
      ("11", "1110001010000010", "0101101111110101", "1111101111110111"), -- i=3551
      ("00", "1010001110110101", "1001011110100101", "0011101101011010"), -- i=3552
      ("01", "1010001110110101", "1001011110100101", "0000110000010000"), -- i=3553
      ("10", "1010001110110101", "1001011110100101", "1000001110100101"), -- i=3554
      ("11", "1010001110110101", "1001011110100101", "1011011110110101"), -- i=3555
      ("00", "1110010011100111", "1100011111010111", "1010110010111110"), -- i=3556
      ("01", "1110010011100111", "1100011111010111", "0001110100010000"), -- i=3557
      ("10", "1110010011100111", "1100011111010111", "1100010011000111"), -- i=3558
      ("11", "1110010011100111", "1100011111010111", "1110011111110111"), -- i=3559
      ("00", "1001110111111100", "1001011000001010", "0011010000000110"), -- i=3560
      ("01", "1001110111111100", "1001011000001010", "0000011111110010"), -- i=3561
      ("10", "1001110111111100", "1001011000001010", "1001010000001000"), -- i=3562
      ("11", "1001110111111100", "1001011000001010", "1001111111111110"), -- i=3563
      ("00", "1110000101010111", "1100100010100001", "1010100111111000"), -- i=3564
      ("01", "1110000101010111", "1100100010100001", "0001100010110110"), -- i=3565
      ("10", "1110000101010111", "1100100010100001", "1100000000000001"), -- i=3566
      ("11", "1110000101010111", "1100100010100001", "1110100111110111"), -- i=3567
      ("00", "1101111001110000", "1011010010011010", "1001001100001010"), -- i=3568
      ("01", "1101111001110000", "1011010010011010", "0010100111010110"), -- i=3569
      ("10", "1101111001110000", "1011010010011010", "1001010000010000"), -- i=3570
      ("11", "1101111001110000", "1011010010011010", "1111111011111010"), -- i=3571
      ("00", "1000100110001111", "0100101111000010", "1101010101010001"), -- i=3572
      ("01", "1000100110001111", "0100101111000010", "0011110111001101"), -- i=3573
      ("10", "1000100110001111", "0100101111000010", "0000100110000010"), -- i=3574
      ("11", "1000100110001111", "0100101111000010", "1100101111001111"), -- i=3575
      ("00", "0101010001010110", "1111110101111100", "0101000111010010"), -- i=3576
      ("01", "0101010001010110", "1111110101111100", "0101011011011010"), -- i=3577
      ("10", "0101010001010110", "1111110101111100", "0101010001010100"), -- i=3578
      ("11", "0101010001010110", "1111110101111100", "1111110101111110"), -- i=3579
      ("00", "1101010011100111", "0000111110100101", "1110010010001100"), -- i=3580
      ("01", "1101010011100111", "0000111110100101", "1100010101000010"), -- i=3581
      ("10", "1101010011100111", "0000111110100101", "0000010010100101"), -- i=3582
      ("11", "1101010011100111", "0000111110100101", "1101111111100111"), -- i=3583
      ("00", "0001110011110000", "0100100000000101", "0110010011110101"), -- i=3584
      ("01", "0001110011110000", "0100100000000101", "1101010011101011"), -- i=3585
      ("10", "0001110011110000", "0100100000000101", "0000100000000000"), -- i=3586
      ("11", "0001110011110000", "0100100000000101", "0101110011110101"), -- i=3587
      ("00", "0001100000001101", "1111100000111101", "0001000001001010"), -- i=3588
      ("01", "0001100000001101", "1111100000111101", "0001111111010000"), -- i=3589
      ("10", "0001100000001101", "1111100000111101", "0001100000001101"), -- i=3590
      ("11", "0001100000001101", "1111100000111101", "1111100000111101"), -- i=3591
      ("00", "1010011010101100", "1111010110111011", "1001110001100111"), -- i=3592
      ("01", "1010011010101100", "1111010110111011", "1011000011110001"), -- i=3593
      ("10", "1010011010101100", "1111010110111011", "1010010010101000"), -- i=3594
      ("11", "1010011010101100", "1111010110111011", "1111011110111111"), -- i=3595
      ("00", "0111100111001100", "0010011111111010", "1010000111000110"), -- i=3596
      ("01", "0111100111001100", "0010011111111010", "0101000111010010"), -- i=3597
      ("10", "0111100111001100", "0010011111111010", "0010000111001000"), -- i=3598
      ("11", "0111100111001100", "0010011111111010", "0111111111111110"), -- i=3599
      ("00", "0111000100001010", "0000000001100111", "0111000101110001"), -- i=3600
      ("01", "0111000100001010", "0000000001100111", "0111000010100011"), -- i=3601
      ("10", "0111000100001010", "0000000001100111", "0000000000000010"), -- i=3602
      ("11", "0111000100001010", "0000000001100111", "0111000101101111"), -- i=3603
      ("00", "0111100101111011", "1111010001010011", "0110110111001110"), -- i=3604
      ("01", "0111100101111011", "1111010001010011", "1000010100101000"), -- i=3605
      ("10", "0111100101111011", "1111010001010011", "0111000001010011"), -- i=3606
      ("11", "0111100101111011", "1111010001010011", "1111110101111011"), -- i=3607
      ("00", "1000110101101011", "0111100100001001", "0000011001110100"), -- i=3608
      ("01", "1000110101101011", "0111100100001001", "0001010001100010"), -- i=3609
      ("10", "1000110101101011", "0111100100001001", "0000100100001001"), -- i=3610
      ("11", "1000110101101011", "0111100100001001", "1111110101101011"), -- i=3611
      ("00", "0111010011110000", "1100100001000110", "0011110100110110"), -- i=3612
      ("01", "0111010011110000", "1100100001000110", "1010110010101010"), -- i=3613
      ("10", "0111010011110000", "1100100001000110", "0100000001000000"), -- i=3614
      ("11", "0111010011110000", "1100100001000110", "1111110011110110"), -- i=3615
      ("00", "1001001001010001", "0000011010111000", "1001100100001001"), -- i=3616
      ("01", "1001001001010001", "0000011010111000", "1000101110011001"), -- i=3617
      ("10", "1001001001010001", "0000011010111000", "0000001000010000"), -- i=3618
      ("11", "1001001001010001", "0000011010111000", "1001011011111001"), -- i=3619
      ("00", "0011110100010001", "0010101010000000", "0110011110010001"), -- i=3620
      ("01", "0011110100010001", "0010101010000000", "0001001010010001"), -- i=3621
      ("10", "0011110100010001", "0010101010000000", "0010100000000000"), -- i=3622
      ("11", "0011110100010001", "0010101010000000", "0011111110010001"), -- i=3623
      ("00", "1010011110111000", "0000101110101011", "1011001101100011"), -- i=3624
      ("01", "1010011110111000", "0000101110101011", "1001110000001101"), -- i=3625
      ("10", "1010011110111000", "0000101110101011", "0000001110101000"), -- i=3626
      ("11", "1010011110111000", "0000101110101011", "1010111110111011"), -- i=3627
      ("00", "1101000101011101", "0110100000011001", "0011100101110110"), -- i=3628
      ("01", "1101000101011101", "0110100000011001", "0110100101000100"), -- i=3629
      ("10", "1101000101011101", "0110100000011001", "0100000000011001"), -- i=3630
      ("11", "1101000101011101", "0110100000011001", "1111100101011101"), -- i=3631
      ("00", "1011000010010000", "1101011000001010", "1000011010011010"), -- i=3632
      ("01", "1011000010010000", "1101011000001010", "1101101010000110"), -- i=3633
      ("10", "1011000010010000", "1101011000001010", "1001000000000000"), -- i=3634
      ("11", "1011000010010000", "1101011000001010", "1111011010011010"), -- i=3635
      ("00", "0100110000000101", "1101100000000010", "0010010000000111"), -- i=3636
      ("01", "0100110000000101", "1101100000000010", "0111010000000011"), -- i=3637
      ("10", "0100110000000101", "1101100000000010", "0100100000000000"), -- i=3638
      ("11", "0100110000000101", "1101100000000010", "1101110000000111"), -- i=3639
      ("00", "0101101010001110", "1010100101000000", "0000001111001110"), -- i=3640
      ("01", "0101101010001110", "1010100101000000", "1011000101001110"), -- i=3641
      ("10", "0101101010001110", "1010100101000000", "0000100000000000"), -- i=3642
      ("11", "0101101010001110", "1010100101000000", "1111101111001110"), -- i=3643
      ("00", "1110000101110000", "0100011010011101", "0010100000001101"), -- i=3644
      ("01", "1110000101110000", "0100011010011101", "1001101011010011"), -- i=3645
      ("10", "1110000101110000", "0100011010011101", "0100000000010000"), -- i=3646
      ("11", "1110000101110000", "0100011010011101", "1110011111111101"), -- i=3647
      ("00", "0000101011001100", "0111101111011100", "1000011010101000"), -- i=3648
      ("01", "0000101011001100", "0111101111011100", "1000111011110000"), -- i=3649
      ("10", "0000101011001100", "0111101111011100", "0000101011001100"), -- i=3650
      ("11", "0000101011001100", "0111101111011100", "0111101111011100"), -- i=3651
      ("00", "1001011101000011", "1101110000100010", "0111001101100101"), -- i=3652
      ("01", "1001011101000011", "1101110000100010", "1011101100100001"), -- i=3653
      ("10", "1001011101000011", "1101110000100010", "1001010000000010"), -- i=3654
      ("11", "1001011101000011", "1101110000100010", "1101111101100011"), -- i=3655
      ("00", "0011001011110001", "1111110101010010", "0011000001000011"), -- i=3656
      ("01", "0011001011110001", "1111110101010010", "0011010110011111"), -- i=3657
      ("10", "0011001011110001", "1111110101010010", "0011000001010000"), -- i=3658
      ("11", "0011001011110001", "1111110101010010", "1111111111110011"), -- i=3659
      ("00", "0000000001001110", "1011101110111000", "1011110000000110"), -- i=3660
      ("01", "0000000001001110", "1011101110111000", "0100010010010110"), -- i=3661
      ("10", "0000000001001110", "1011101110111000", "0000000000001000"), -- i=3662
      ("11", "0000000001001110", "1011101110111000", "1011101111111110"), -- i=3663
      ("00", "1001011111100010", "1101011000100000", "0110111000000010"), -- i=3664
      ("01", "1001011111100010", "1101011000100000", "1100000111000010"), -- i=3665
      ("10", "1001011111100010", "1101011000100000", "1001011000100000"), -- i=3666
      ("11", "1001011111100010", "1101011000100000", "1101011111100010"), -- i=3667
      ("00", "1101101111101111", "1010110001110100", "1000100001100011"), -- i=3668
      ("01", "1101101111101111", "1010110001110100", "0010111101111011"), -- i=3669
      ("10", "1101101111101111", "1010110001110100", "1000100001100100"), -- i=3670
      ("11", "1101101111101111", "1010110001110100", "1111111111111111"), -- i=3671
      ("00", "0111100000110000", "0001110000011011", "1001010001001011"), -- i=3672
      ("01", "0111100000110000", "0001110000011011", "0101110000010101"), -- i=3673
      ("10", "0111100000110000", "0001110000011011", "0001100000010000"), -- i=3674
      ("11", "0111100000110000", "0001110000011011", "0111110000111011"), -- i=3675
      ("00", "1111000011000010", "0101100010100011", "0100100101100101"), -- i=3676
      ("01", "1111000011000010", "0101100010100011", "1001100000011111"), -- i=3677
      ("10", "1111000011000010", "0101100010100011", "0101000010000010"), -- i=3678
      ("11", "1111000011000010", "0101100010100011", "1111100011100011"), -- i=3679
      ("00", "0100110110111000", "1010001111111101", "1111000110110101"), -- i=3680
      ("01", "0100110110111000", "1010001111111101", "1010100110111011"), -- i=3681
      ("10", "0100110110111000", "1010001111111101", "0000000110111000"), -- i=3682
      ("11", "0100110110111000", "1010001111111101", "1110111111111101"), -- i=3683
      ("00", "1101101111001001", "0001001100000110", "1110111011001111"), -- i=3684
      ("01", "1101101111001001", "0001001100000110", "1100100011000011"), -- i=3685
      ("10", "1101101111001001", "0001001100000110", "0001001100000000"), -- i=3686
      ("11", "1101101111001001", "0001001100000110", "1101101111001111"), -- i=3687
      ("00", "0001101101000011", "0011000001110100", "0100101110110111"), -- i=3688
      ("01", "0001101101000011", "0011000001110100", "1110101011001111"), -- i=3689
      ("10", "0001101101000011", "0011000001110100", "0001000001000000"), -- i=3690
      ("11", "0001101101000011", "0011000001110100", "0011101101110111"), -- i=3691
      ("00", "1101011001011000", "1001110011110101", "0111001101001101"), -- i=3692
      ("01", "1101011001011000", "1001110011110101", "0011100101100011"), -- i=3693
      ("10", "1101011001011000", "1001110011110101", "1001010001010000"), -- i=3694
      ("11", "1101011001011000", "1001110011110101", "1101111011111101"), -- i=3695
      ("00", "1101010000000000", "0111111000111001", "0101001000111001"), -- i=3696
      ("01", "1101010000000000", "0111111000111001", "0101010111000111"), -- i=3697
      ("10", "1101010000000000", "0111111000111001", "0101010000000000"), -- i=3698
      ("11", "1101010000000000", "0111111000111001", "1111111000111001"), -- i=3699
      ("00", "1010011001011011", "0001101110000101", "1100000111100000"), -- i=3700
      ("01", "1010011001011011", "0001101110000101", "1000101011010110"), -- i=3701
      ("10", "1010011001011011", "0001101110000101", "0000001000000001"), -- i=3702
      ("11", "1010011001011011", "0001101110000101", "1011111111011111"), -- i=3703
      ("00", "0111000000110111", "1101010000000101", "0100010000111100"), -- i=3704
      ("01", "0111000000110111", "1101010000000101", "1001110000110010"), -- i=3705
      ("10", "0111000000110111", "1101010000000101", "0101000000000101"), -- i=3706
      ("11", "0111000000110111", "1101010000000101", "1111010000110111"), -- i=3707
      ("00", "0000010111100010", "0100010100100101", "0100101100000111"), -- i=3708
      ("01", "0000010111100010", "0100010100100101", "1100000010111101"), -- i=3709
      ("10", "0000010111100010", "0100010100100101", "0000010100100000"), -- i=3710
      ("11", "0000010111100010", "0100010100100101", "0100010111100111"), -- i=3711
      ("00", "1010111110001101", "0000110001100010", "1011101111101111"), -- i=3712
      ("01", "1010111110001101", "0000110001100010", "1010001100101011"), -- i=3713
      ("10", "1010111110001101", "0000110001100010", "0000110000000000"), -- i=3714
      ("11", "1010111110001101", "0000110001100010", "1010111111101111"), -- i=3715
      ("00", "1100111111111011", "1101010001011001", "1010010001010100"), -- i=3716
      ("01", "1100111111111011", "1101010001011001", "1111101110100010"), -- i=3717
      ("10", "1100111111111011", "1101010001011001", "1100010001011001"), -- i=3718
      ("11", "1100111111111011", "1101010001011001", "1101111111111011"), -- i=3719
      ("00", "0101111010101111", "0000011010100100", "0110010101010011"), -- i=3720
      ("01", "0101111010101111", "0000011010100100", "0101100000001011"), -- i=3721
      ("10", "0101111010101111", "0000011010100100", "0000011010100100"), -- i=3722
      ("11", "0101111010101111", "0000011010100100", "0101111010101111"), -- i=3723
      ("00", "0010101001000000", "0111011101111010", "1010000110111010"), -- i=3724
      ("01", "0010101001000000", "0111011101111010", "1011001011000110"), -- i=3725
      ("10", "0010101001000000", "0111011101111010", "0010001001000000"), -- i=3726
      ("11", "0010101001000000", "0111011101111010", "0111111101111010"), -- i=3727
      ("00", "0011001101000101", "0000101110100010", "0011111011100111"), -- i=3728
      ("01", "0011001101000101", "0000101110100010", "0010011110100011"), -- i=3729
      ("10", "0011001101000101", "0000101110100010", "0000001100000000"), -- i=3730
      ("11", "0011001101000101", "0000101110100010", "0011101111100111"), -- i=3731
      ("00", "1011001110101001", "1100100010101111", "0111110001011000"), -- i=3732
      ("01", "1011001110101001", "1100100010101111", "1110101011111010"), -- i=3733
      ("10", "1011001110101001", "1100100010101111", "1000000010101001"), -- i=3734
      ("11", "1011001110101001", "1100100010101111", "1111101110101111"), -- i=3735
      ("00", "1111011001111100", "1111100111100010", "1111000001011110"), -- i=3736
      ("01", "1111011001111100", "1111100111100010", "1111110010011010"), -- i=3737
      ("10", "1111011001111100", "1111100111100010", "1111000001100000"), -- i=3738
      ("11", "1111011001111100", "1111100111100010", "1111111111111110"), -- i=3739
      ("00", "0111101010000111", "0101010001110110", "1100111011111101"), -- i=3740
      ("01", "0111101010000111", "0101010001110110", "0010011000010001"), -- i=3741
      ("10", "0111101010000111", "0101010001110110", "0101000000000110"), -- i=3742
      ("11", "0111101010000111", "0101010001110110", "0111111011110111"), -- i=3743
      ("00", "1100001110011001", "1111110001010001", "1011111111101010"), -- i=3744
      ("01", "1100001110011001", "1111110001010001", "1100011101001000"), -- i=3745
      ("10", "1100001110011001", "1111110001010001", "1100000000010001"), -- i=3746
      ("11", "1100001110011001", "1111110001010001", "1111111111011001"), -- i=3747
      ("00", "0001110010111000", "0101100001111111", "0111010100110111"), -- i=3748
      ("01", "0001110010111000", "0101100001111111", "1100010000111001"), -- i=3749
      ("10", "0001110010111000", "0101100001111111", "0001100000111000"), -- i=3750
      ("11", "0001110010111000", "0101100001111111", "0101110011111111"), -- i=3751
      ("00", "1001010101000110", "0010010111010101", "1011101100011011"), -- i=3752
      ("01", "1001010101000110", "0010010111010101", "0110111101110001"), -- i=3753
      ("10", "1001010101000110", "0010010111010101", "0000010101000100"), -- i=3754
      ("11", "1001010101000110", "0010010111010101", "1011010111010111"), -- i=3755
      ("00", "1111111001110101", "1010111110101110", "1010111000100011"), -- i=3756
      ("01", "1111111001110101", "1010111110101110", "0100111011000111"), -- i=3757
      ("10", "1111111001110101", "1010111110101110", "1010111000100100"), -- i=3758
      ("11", "1111111001110101", "1010111110101110", "1111111111111111"), -- i=3759
      ("00", "0011100110100010", "1000101100110000", "1100010011010010"), -- i=3760
      ("01", "0011100110100010", "1000101100110000", "1010111001110010"), -- i=3761
      ("10", "0011100110100010", "1000101100110000", "0000100100100000"), -- i=3762
      ("11", "0011100110100010", "1000101100110000", "1011101110110010"), -- i=3763
      ("00", "1111010101010000", "0101001101111011", "0100100011001011"), -- i=3764
      ("01", "1111010101010000", "0101001101111011", "1010000111010101"), -- i=3765
      ("10", "1111010101010000", "0101001101111011", "0101000101010000"), -- i=3766
      ("11", "1111010101010000", "0101001101111011", "1111011101111011"), -- i=3767
      ("00", "0000101001000111", "0101110000010011", "0110011001011010"), -- i=3768
      ("01", "0000101001000111", "0101110000010011", "1010111000110100"), -- i=3769
      ("10", "0000101001000111", "0101110000010011", "0000100000000011"), -- i=3770
      ("11", "0000101001000111", "0101110000010011", "0101111001010111"), -- i=3771
      ("00", "0001111000111101", "1111011000011000", "0001010001010101"), -- i=3772
      ("01", "0001111000111101", "1111011000011000", "0010100000100101"), -- i=3773
      ("10", "0001111000111101", "1111011000011000", "0001011000011000"), -- i=3774
      ("11", "0001111000111101", "1111011000011000", "1111111000111101"), -- i=3775
      ("00", "0111001010111110", "0000101101100000", "0111111000011110"), -- i=3776
      ("01", "0111001010111110", "0000101101100000", "0110011101011110"), -- i=3777
      ("10", "0111001010111110", "0000101101100000", "0000001000100000"), -- i=3778
      ("11", "0111001010111110", "0000101101100000", "0111101111111110"), -- i=3779
      ("00", "1101011011000011", "0111101111111101", "0101001011000000"), -- i=3780
      ("01", "1101011011000011", "0111101111111101", "0101101011000110"), -- i=3781
      ("10", "1101011011000011", "0111101111111101", "0101001011000001"), -- i=3782
      ("11", "1101011011000011", "0111101111111101", "1111111111111111"), -- i=3783
      ("00", "0110010100100000", "1100110111011111", "0011001011111111"), -- i=3784
      ("01", "0110010100100000", "1100110111011111", "1001011101000001"), -- i=3785
      ("10", "0110010100100000", "1100110111011111", "0100010100000000"), -- i=3786
      ("11", "0110010100100000", "1100110111011111", "1110110111111111"), -- i=3787
      ("00", "1111101010100110", "1000011011010100", "1000000101111010"), -- i=3788
      ("01", "1111101010100110", "1000011011010100", "0111001111010010"), -- i=3789
      ("10", "1111101010100110", "1000011011010100", "1000001010000100"), -- i=3790
      ("11", "1111101010100110", "1000011011010100", "1111111011110110"), -- i=3791
      ("00", "0101100111010111", "1001011000001001", "1110111111100000"), -- i=3792
      ("01", "0101100111010111", "1001011000001001", "1100001111001110"), -- i=3793
      ("10", "0101100111010111", "1001011000001001", "0001000000000001"), -- i=3794
      ("11", "0101100111010111", "1001011000001001", "1101111111011111"), -- i=3795
      ("00", "1001100010110110", "1101011011100011", "0110111110011001"), -- i=3796
      ("01", "1001100010110110", "1101011011100011", "1100000111010011"), -- i=3797
      ("10", "1001100010110110", "1101011011100011", "1001000010100010"), -- i=3798
      ("11", "1001100010110110", "1101011011100011", "1101111011110111"), -- i=3799
      ("00", "0101110011000000", "0011101010001011", "1001011101001011"), -- i=3800
      ("01", "0101110011000000", "0011101010001011", "0010001000110101"), -- i=3801
      ("10", "0101110011000000", "0011101010001011", "0001100010000000"), -- i=3802
      ("11", "0101110011000000", "0011101010001011", "0111111011001011"), -- i=3803
      ("00", "0100101001111111", "0000001101011111", "0100110111011110"), -- i=3804
      ("01", "0100101001111111", "0000001101011111", "0100011100100000"), -- i=3805
      ("10", "0100101001111111", "0000001101011111", "0000001001011111"), -- i=3806
      ("11", "0100101001111111", "0000001101011111", "0100101101111111"), -- i=3807
      ("00", "1111011100101001", "1010010010111000", "1001101111100001"), -- i=3808
      ("01", "1111011100101001", "1010010010111000", "0101001001110001"), -- i=3809
      ("10", "1111011100101001", "1010010010111000", "1010010000101000"), -- i=3810
      ("11", "1111011100101001", "1010010010111000", "1111011110111001"), -- i=3811
      ("00", "0011110000011101", "1110110101011111", "0010100101111100"), -- i=3812
      ("01", "0011110000011101", "1110110101011111", "0100111010111110"), -- i=3813
      ("10", "0011110000011101", "1110110101011111", "0010110000011101"), -- i=3814
      ("11", "0011110000011101", "1110110101011111", "1111110101011111"), -- i=3815
      ("00", "0111101101011001", "1011101100001101", "0011011001100110"), -- i=3816
      ("01", "0111101101011001", "1011101100001101", "1100000001001100"), -- i=3817
      ("10", "0111101101011001", "1011101100001101", "0011101100001001"), -- i=3818
      ("11", "0111101101011001", "1011101100001101", "1111101101011101"), -- i=3819
      ("00", "1011101001100010", "0101110001000000", "0001011010100010"), -- i=3820
      ("01", "1011101001100010", "0101110001000000", "0101111000100010"), -- i=3821
      ("10", "1011101001100010", "0101110001000000", "0001100001000000"), -- i=3822
      ("11", "1011101001100010", "0101110001000000", "1111111001100010"), -- i=3823
      ("00", "0101001110101101", "0011101101101110", "1000111100011011"), -- i=3824
      ("01", "0101001110101101", "0011101101101110", "0001100000111111"), -- i=3825
      ("10", "0101001110101101", "0011101101101110", "0001001100101100"), -- i=3826
      ("11", "0101001110101101", "0011101101101110", "0111101111101111"), -- i=3827
      ("00", "1100111100001100", "0110010111000000", "0011010011001100"), -- i=3828
      ("01", "1100111100001100", "0110010111000000", "0110100101001100"), -- i=3829
      ("10", "1100111100001100", "0110010111000000", "0100010100000000"), -- i=3830
      ("11", "1100111100001100", "0110010111000000", "1110111111001100"), -- i=3831
      ("00", "0111110001110011", "1101111111001110", "0101110001000001"), -- i=3832
      ("01", "0111110001110011", "1101111111001110", "1001110010100101"), -- i=3833
      ("10", "0111110001110011", "1101111111001110", "0101110001000010"), -- i=3834
      ("11", "0111110001110011", "1101111111001110", "1111111111111111"), -- i=3835
      ("00", "0000101111010001", "1001111100100110", "1010101011110111"), -- i=3836
      ("01", "0000101111010001", "1001111100100110", "0110110010101011"), -- i=3837
      ("10", "0000101111010001", "1001111100100110", "0000101100000000"), -- i=3838
      ("11", "0000101111010001", "1001111100100110", "1001111111110111"), -- i=3839
      ("00", "0011110100001101", "1111011101100101", "0011010001110010"), -- i=3840
      ("01", "0011110100001101", "1111011101100101", "0100010110101000"), -- i=3841
      ("10", "0011110100001101", "1111011101100101", "0011010100000101"), -- i=3842
      ("11", "0011110100001101", "1111011101100101", "1111111101101101"), -- i=3843
      ("00", "0010011001011110", "1001100000100111", "1011111010000101"), -- i=3844
      ("01", "0010011001011110", "1001100000100111", "1000111000110111"), -- i=3845
      ("10", "0010011001011110", "1001100000100111", "0000000000000110"), -- i=3846
      ("11", "0010011001011110", "1001100000100111", "1011111001111111"), -- i=3847
      ("00", "1000101000001010", "0001010110100011", "1001111110101101"), -- i=3848
      ("01", "1000101000001010", "0001010110100011", "0111010001100111"), -- i=3849
      ("10", "1000101000001010", "0001010110100011", "0000000000000010"), -- i=3850
      ("11", "1000101000001010", "0001010110100011", "1001111110101011"), -- i=3851
      ("00", "0111000010101000", "1100101101111011", "0011110000100011"), -- i=3852
      ("01", "0111000010101000", "1100101101111011", "1010010100101101"), -- i=3853
      ("10", "0111000010101000", "1100101101111011", "0100000000101000"), -- i=3854
      ("11", "0111000010101000", "1100101101111011", "1111101111111011"), -- i=3855
      ("00", "0011011100110010", "1001011110000111", "1100111010111001"), -- i=3856
      ("01", "0011011100110010", "1001011110000111", "1001111110101011"), -- i=3857
      ("10", "0011011100110010", "1001011110000111", "0001011100000010"), -- i=3858
      ("11", "0011011100110010", "1001011110000111", "1011011110110111"), -- i=3859
      ("00", "1000101000101010", "0000010000110111", "1000111001100001"), -- i=3860
      ("01", "1000101000101010", "0000010000110111", "1000010111110011"), -- i=3861
      ("10", "1000101000101010", "0000010000110111", "0000000000100010"), -- i=3862
      ("11", "1000101000101010", "0000010000110111", "1000111000111111"), -- i=3863
      ("00", "0100010111000101", "1000011100000011", "1100110011001000"), -- i=3864
      ("01", "0100010111000101", "1000011100000011", "1011111011000010"), -- i=3865
      ("10", "0100010111000101", "1000011100000011", "0000010100000001"), -- i=3866
      ("11", "0100010111000101", "1000011100000011", "1100011111000111"), -- i=3867
      ("00", "1101111111011011", "0011001001101110", "0001001001001001"), -- i=3868
      ("01", "1101111111011011", "0011001001101110", "1010110101101101"), -- i=3869
      ("10", "1101111111011011", "0011001001101110", "0001001001001010"), -- i=3870
      ("11", "1101111111011011", "0011001001101110", "1111111111111111"), -- i=3871
      ("00", "0010100001100000", "1101001110011100", "1111101111111100"), -- i=3872
      ("01", "0010100001100000", "1101001110011100", "0101010011000100"), -- i=3873
      ("10", "0010100001100000", "1101001110011100", "0000000000000000"), -- i=3874
      ("11", "0010100001100000", "1101001110011100", "1111101111111100"), -- i=3875
      ("00", "1011001000010001", "1100110010110100", "0111111011000101"), -- i=3876
      ("01", "1011001000010001", "1100110010110100", "1110010101011101"), -- i=3877
      ("10", "1011001000010001", "1100110010110100", "1000000000010000"), -- i=3878
      ("11", "1011001000010001", "1100110010110100", "1111111010110101"), -- i=3879
      ("00", "1100101101000010", "1110111001101011", "1011100110101101"), -- i=3880
      ("01", "1100101101000010", "1110111001101011", "1101110011010111"), -- i=3881
      ("10", "1100101101000010", "1110111001101011", "1100101001000010"), -- i=3882
      ("11", "1100101101000010", "1110111001101011", "1110111101101011"), -- i=3883
      ("00", "0110000010001110", "0010011101101101", "1000011111111011"), -- i=3884
      ("01", "0110000010001110", "0010011101101101", "0011100100100001"), -- i=3885
      ("10", "0110000010001110", "0010011101101101", "0010000000001100"), -- i=3886
      ("11", "0110000010001110", "0010011101101101", "0110011111101111"), -- i=3887
      ("00", "1000110011101111", "1001011100101010", "0010010000011001"), -- i=3888
      ("01", "1000110011101111", "1001011100101010", "1111010111000101"), -- i=3889
      ("10", "1000110011101111", "1001011100101010", "1000010000101010"), -- i=3890
      ("11", "1000110011101111", "1001011100101010", "1001111111101111"), -- i=3891
      ("00", "1010111001100010", "1001111000011100", "0100110001111110"), -- i=3892
      ("01", "1010111001100010", "1001111000011100", "0001000001000110"), -- i=3893
      ("10", "1010111001100010", "1001111000011100", "1000111000000000"), -- i=3894
      ("11", "1010111001100010", "1001111000011100", "1011111001111110"), -- i=3895
      ("00", "0001100001101111", "0000111011111010", "0010011101101001"), -- i=3896
      ("01", "0001100001101111", "0000111011111010", "0000100101110101"), -- i=3897
      ("10", "0001100001101111", "0000111011111010", "0000100001101010"), -- i=3898
      ("11", "0001100001101111", "0000111011111010", "0001111011111111"), -- i=3899
      ("00", "1000100010000000", "0000011000010010", "1000111010010010"), -- i=3900
      ("01", "1000100010000000", "0000011000010010", "1000001001101110"), -- i=3901
      ("10", "1000100010000000", "0000011000010010", "0000000000000000"), -- i=3902
      ("11", "1000100010000000", "0000011000010010", "1000111010010010"), -- i=3903
      ("00", "0011111110010000", "1111010100001000", "0011010010011000"), -- i=3904
      ("01", "0011111110010000", "1111010100001000", "0100101010001000"), -- i=3905
      ("10", "0011111110010000", "1111010100001000", "0011010100000000"), -- i=3906
      ("11", "0011111110010000", "1111010100001000", "1111111110011000"), -- i=3907
      ("00", "1001101100001011", "1010010100101100", "0100000000110111"), -- i=3908
      ("01", "1001101100001011", "1010010100101100", "1111010111011111"), -- i=3909
      ("10", "1001101100001011", "1010010100101100", "1000000100001000"), -- i=3910
      ("11", "1001101100001011", "1010010100101100", "1011111100101111"), -- i=3911
      ("00", "1000100100000001", "1100100000111110", "0101000100111111"), -- i=3912
      ("01", "1000100100000001", "1100100000111110", "1100000011000011"), -- i=3913
      ("10", "1000100100000001", "1100100000111110", "1000100000000000"), -- i=3914
      ("11", "1000100100000001", "1100100000111110", "1100100100111111"), -- i=3915
      ("00", "1010101011001110", "1101001010001001", "0111110101010111"), -- i=3916
      ("01", "1010101011001110", "1101001010001001", "1101100001000101"), -- i=3917
      ("10", "1010101011001110", "1101001010001001", "1000001010001000"), -- i=3918
      ("11", "1010101011001110", "1101001010001001", "1111101011001111"), -- i=3919
      ("00", "0010001100100111", "0110100010100111", "1000101111001110"), -- i=3920
      ("01", "0010001100100111", "0110100010100111", "1011101010000000"), -- i=3921
      ("10", "0010001100100111", "0110100010100111", "0010000000100111"), -- i=3922
      ("11", "0010001100100111", "0110100010100111", "0110101110100111"), -- i=3923
      ("00", "0011100101100100", "0111101001100001", "1011001111000101"), -- i=3924
      ("01", "0011100101100100", "0111101001100001", "1011111100000011"), -- i=3925
      ("10", "0011100101100100", "0111101001100001", "0011100001100000"), -- i=3926
      ("11", "0011100101100100", "0111101001100001", "0111101101100101"), -- i=3927
      ("00", "0101000111110110", "1111101000110111", "0100110000101101"), -- i=3928
      ("01", "0101000111110110", "1111101000110111", "0101011110111111"), -- i=3929
      ("10", "0101000111110110", "1111101000110111", "0101000000110110"), -- i=3930
      ("11", "0101000111110110", "1111101000110111", "1111101111110111"), -- i=3931
      ("00", "0111001111111101", "1111100101101000", "0110110101100101"), -- i=3932
      ("01", "0111001111111101", "1111100101101000", "0111101010010101"), -- i=3933
      ("10", "0111001111111101", "1111100101101000", "0111000101101000"), -- i=3934
      ("11", "0111001111111101", "1111100101101000", "1111101111111101"), -- i=3935
      ("00", "0011101100111111", "0011101000010000", "0111010101001111"), -- i=3936
      ("01", "0011101100111111", "0011101000010000", "0000000100101111"), -- i=3937
      ("10", "0011101100111111", "0011101000010000", "0011101000010000"), -- i=3938
      ("11", "0011101100111111", "0011101000010000", "0011101100111111"), -- i=3939
      ("00", "1100110111001000", "0010011101100111", "1111010100101111"), -- i=3940
      ("01", "1100110111001000", "0010011101100111", "1010011001100001"), -- i=3941
      ("10", "1100110111001000", "0010011101100111", "0000010101000000"), -- i=3942
      ("11", "1100110111001000", "0010011101100111", "1110111111101111"), -- i=3943
      ("00", "0010101000110010", "1010111010001101", "1101100010111111"), -- i=3944
      ("01", "0010101000110010", "1010111010001101", "0111101110100101"), -- i=3945
      ("10", "0010101000110010", "1010111010001101", "0010101000000000"), -- i=3946
      ("11", "0010101000110010", "1010111010001101", "1010111010111111"), -- i=3947
      ("00", "1111000001101001", "1111001111110111", "1110010001100000"), -- i=3948
      ("01", "1111000001101001", "1111001111110111", "1111110001110010"), -- i=3949
      ("10", "1111000001101001", "1111001111110111", "1111000001100001"), -- i=3950
      ("11", "1111000001101001", "1111001111110111", "1111001111111111"), -- i=3951
      ("00", "0000000000001011", "0001100110010010", "0001100110011101"), -- i=3952
      ("01", "0000000000001011", "0001100110010010", "1110011001111001"), -- i=3953
      ("10", "0000000000001011", "0001100110010010", "0000000000000010"), -- i=3954
      ("11", "0000000000001011", "0001100110010010", "0001100110011011"), -- i=3955
      ("00", "1101111000001101", "1010101110000000", "1000100110001101"), -- i=3956
      ("01", "1101111000001101", "1010101110000000", "0011001010001101"), -- i=3957
      ("10", "1101111000001101", "1010101110000000", "1000101000000000"), -- i=3958
      ("11", "1101111000001101", "1010101110000000", "1111111110001101"), -- i=3959
      ("00", "1000110100101001", "0011101111111011", "1100100100100100"), -- i=3960
      ("01", "1000110100101001", "0011101111111011", "0101000100101110"), -- i=3961
      ("10", "1000110100101001", "0011101111111011", "0000100100101001"), -- i=3962
      ("11", "1000110100101001", "0011101111111011", "1011111111111011"), -- i=3963
      ("00", "0011100111111101", "1101010111110010", "0000111111101111"), -- i=3964
      ("01", "0011100111111101", "1101010111110010", "0110010000001011"), -- i=3965
      ("10", "0011100111111101", "1101010111110010", "0001000111110000"), -- i=3966
      ("11", "0011100111111101", "1101010111110010", "1111110111111111"), -- i=3967
      ("00", "1111101011111111", "0100100000100111", "0100001100100110"), -- i=3968
      ("01", "1111101011111111", "0100100000100111", "1011001011011000"), -- i=3969
      ("10", "1111101011111111", "0100100000100111", "0100100000100111"), -- i=3970
      ("11", "1111101011111111", "0100100000100111", "1111101011111111"), -- i=3971
      ("00", "1010110111000011", "1010001111011010", "0101000110011101"), -- i=3972
      ("01", "1010110111000011", "1010001111011010", "0000100111101001"), -- i=3973
      ("10", "1010110111000011", "1010001111011010", "1010000111000010"), -- i=3974
      ("11", "1010110111000011", "1010001111011010", "1010111111011011"), -- i=3975
      ("00", "0100010010100100", "0101100011101101", "1001110110010001"), -- i=3976
      ("01", "0100010010100100", "0101100011101101", "1110101110110111"), -- i=3977
      ("10", "0100010010100100", "0101100011101101", "0100000010100100"), -- i=3978
      ("11", "0100010010100100", "0101100011101101", "0101110011101101"), -- i=3979
      ("00", "0100101000111111", "0000100110111011", "0101001111111010"), -- i=3980
      ("01", "0100101000111111", "0000100110111011", "0100000010000100"), -- i=3981
      ("10", "0100101000111111", "0000100110111011", "0000100000111011"), -- i=3982
      ("11", "0100101000111111", "0000100110111011", "0100101110111111"), -- i=3983
      ("00", "1111100011111010", "1110000110001100", "1101101010000110"), -- i=3984
      ("01", "1111100011111010", "1110000110001100", "0001011101101110"), -- i=3985
      ("10", "1111100011111010", "1110000110001100", "1110000010001000"), -- i=3986
      ("11", "1111100011111010", "1110000110001100", "1111100111111110"), -- i=3987
      ("00", "1001010101001100", "1111110011100001", "1001001000101101"), -- i=3988
      ("01", "1001010101001100", "1111110011100001", "1001100001101011"), -- i=3989
      ("10", "1001010101001100", "1111110011100001", "1001010001000000"), -- i=3990
      ("11", "1001010101001100", "1111110011100001", "1111110111101101"), -- i=3991
      ("00", "0010011010010111", "0101001001010001", "0111100011101000"), -- i=3992
      ("01", "0010011010010111", "0101001001010001", "1101010001000110"), -- i=3993
      ("10", "0010011010010111", "0101001001010001", "0000001000010001"), -- i=3994
      ("11", "0010011010010111", "0101001001010001", "0111011011010111"), -- i=3995
      ("00", "1010110110111000", "1100000000000100", "0110110110111100"), -- i=3996
      ("01", "1010110110111000", "1100000000000100", "1110110110110100"), -- i=3997
      ("10", "1010110110111000", "1100000000000100", "1000000000000000"), -- i=3998
      ("11", "1010110110111000", "1100000000000100", "1110110110111100"), -- i=3999
      ("00", "0101111100001001", "0001110100001110", "0111110000010111"), -- i=4000
      ("01", "0101111100001001", "0001110100001110", "0100000111111011"), -- i=4001
      ("10", "0101111100001001", "0001110100001110", "0001110100001000"), -- i=4002
      ("11", "0101111100001001", "0001110100001110", "0101111100001111"), -- i=4003
      ("00", "1001000011001110", "1101000101111101", "0110001001001011"), -- i=4004
      ("01", "1001000011001110", "1101000101111101", "1011111101010001"), -- i=4005
      ("10", "1001000011001110", "1101000101111101", "1001000001001100"), -- i=4006
      ("11", "1001000011001110", "1101000101111101", "1101000111111111"), -- i=4007
      ("00", "0011010000001000", "1101101110011111", "0000111110100111"), -- i=4008
      ("01", "0011010000001000", "1101101110011111", "0101100001101001"), -- i=4009
      ("10", "0011010000001000", "1101101110011111", "0001000000001000"), -- i=4010
      ("11", "0011010000001000", "1101101110011111", "1111111110011111"), -- i=4011
      ("00", "0001010110100111", "1101011111100100", "1110110110001011"), -- i=4012
      ("01", "0001010110100111", "1101011111100100", "0011110111000011"), -- i=4013
      ("10", "0001010110100111", "1101011111100100", "0001010110100100"), -- i=4014
      ("11", "0001010110100111", "1101011111100100", "1101011111100111"), -- i=4015
      ("00", "0110111010110111", "1001101000001100", "0000100011000011"), -- i=4016
      ("01", "0110111010110111", "1001101000001100", "1101010010101011"), -- i=4017
      ("10", "0110111010110111", "1001101000001100", "0000101000000100"), -- i=4018
      ("11", "0110111010110111", "1001101000001100", "1111111010111111"), -- i=4019
      ("00", "1010001111110010", "1101110101001001", "1000000100111011"), -- i=4020
      ("01", "1010001111110010", "1101110101001001", "1100011010101001"), -- i=4021
      ("10", "1010001111110010", "1101110101001001", "1000000101000000"), -- i=4022
      ("11", "1010001111110010", "1101110101001001", "1111111111111011"), -- i=4023
      ("00", "1000011000001110", "0010110100010100", "1011001100100010"), -- i=4024
      ("01", "1000011000001110", "0010110100010100", "0101100011111010"), -- i=4025
      ("10", "1000011000001110", "0010110100010100", "0000010000000100"), -- i=4026
      ("11", "1000011000001110", "0010110100010100", "1010111100011110"), -- i=4027
      ("00", "0000010100001100", "0100010001101111", "0100100101111011"), -- i=4028
      ("01", "0000010100001100", "0100010001101111", "1100000010011101"), -- i=4029
      ("10", "0000010100001100", "0100010001101111", "0000010000001100"), -- i=4030
      ("11", "0000010100001100", "0100010001101111", "0100010101101111"), -- i=4031
      ("00", "1000011011111001", "0000110100100111", "1001010000100000"), -- i=4032
      ("01", "1000011011111001", "0000110100100111", "0111100111010010"), -- i=4033
      ("10", "1000011011111001", "0000110100100111", "0000010000100001"), -- i=4034
      ("11", "1000011011111001", "0000110100100111", "1000111111111111"), -- i=4035
      ("00", "1110111101110100", "0010011010111011", "0001011000101111"), -- i=4036
      ("01", "1110111101110100", "0010011010111011", "1100100010111001"), -- i=4037
      ("10", "1110111101110100", "0010011010111011", "0010011000110000"), -- i=4038
      ("11", "1110111101110100", "0010011010111011", "1110111111111111"), -- i=4039
      ("00", "1011010111100100", "0110010100011100", "0001101100000000"), -- i=4040
      ("01", "1011010111100100", "0110010100011100", "0101000011001000"), -- i=4041
      ("10", "1011010111100100", "0110010100011100", "0010010100000100"), -- i=4042
      ("11", "1011010111100100", "0110010100011100", "1111010111111100"), -- i=4043
      ("00", "0001011000001000", "0011010010110010", "0100101010111010"), -- i=4044
      ("01", "0001011000001000", "0011010010110010", "1110000101010110"), -- i=4045
      ("10", "0001011000001000", "0011010010110010", "0001010000000000"), -- i=4046
      ("11", "0001011000001000", "0011010010110010", "0011011010111010"), -- i=4047
      ("00", "1010111010100101", "1110001100101101", "1001000111010010"), -- i=4048
      ("01", "1010111010100101", "1110001100101101", "1100101101111000"), -- i=4049
      ("10", "1010111010100101", "1110001100101101", "1010001000100101"), -- i=4050
      ("11", "1010111010100101", "1110001100101101", "1110111110101101"), -- i=4051
      ("00", "1001010110010011", "1100011001000001", "0101101111010100"), -- i=4052
      ("01", "1001010110010011", "1100011001000001", "1100111101010010"), -- i=4053
      ("10", "1001010110010011", "1100011001000001", "1000010000000001"), -- i=4054
      ("11", "1001010110010011", "1100011001000001", "1101011111010011"), -- i=4055
      ("00", "1010110100001101", "0110000111111011", "0000111100001000"), -- i=4056
      ("01", "1010110100001101", "0110000111111011", "0100101100010010"), -- i=4057
      ("10", "1010110100001101", "0110000111111011", "0010000100001001"), -- i=4058
      ("11", "1010110100001101", "0110000111111011", "1110110111111111"), -- i=4059
      ("00", "1001010010010010", "1000001100101101", "0001011110111111"), -- i=4060
      ("01", "1001010010010010", "1000001100101101", "0001000101100101"), -- i=4061
      ("10", "1001010010010010", "1000001100101101", "1000000000000000"), -- i=4062
      ("11", "1001010010010010", "1000001100101101", "1001011110111111"), -- i=4063
      ("00", "1111010110000111", "1010111010110110", "1010010000111101"), -- i=4064
      ("01", "1111010110000111", "1010111010110110", "0100011011010001"), -- i=4065
      ("10", "1111010110000111", "1010111010110110", "1010010010000110"), -- i=4066
      ("11", "1111010110000111", "1010111010110110", "1111111110110111"), -- i=4067
      ("00", "1100101001001001", "1110111101010110", "1011100110011111"), -- i=4068
      ("01", "1100101001001001", "1110111101010110", "1101101011110011"), -- i=4069
      ("10", "1100101001001001", "1110111101010110", "1100101001000000"), -- i=4070
      ("11", "1100101001001001", "1110111101010110", "1110111101011111"), -- i=4071
      ("00", "0000101010010010", "1000100010011110", "1001001100110000"), -- i=4072
      ("01", "0000101010010010", "1000100010011110", "1000000111110100"), -- i=4073
      ("10", "0000101010010010", "1000100010011110", "0000100010010010"), -- i=4074
      ("11", "0000101010010010", "1000100010011110", "1000101010011110"), -- i=4075
      ("00", "0110101101111001", "0011000110111111", "1001110100111000"), -- i=4076
      ("01", "0110101101111001", "0011000110111111", "0011100110111010"), -- i=4077
      ("10", "0110101101111001", "0011000110111111", "0010000100111001"), -- i=4078
      ("11", "0110101101111001", "0011000110111111", "0111101111111111"), -- i=4079
      ("00", "0111100100000001", "0111010101110100", "1110111001110101"), -- i=4080
      ("01", "0111100100000001", "0111010101110100", "0000001110001101"), -- i=4081
      ("10", "0111100100000001", "0111010101110100", "0111000100000000"), -- i=4082
      ("11", "0111100100000001", "0111010101110100", "0111110101110101"), -- i=4083
      ("00", "1010110001011101", "1010000010000001", "0100110011011110"), -- i=4084
      ("01", "1010110001011101", "1010000010000001", "0000101111011100"), -- i=4085
      ("10", "1010110001011101", "1010000010000001", "1010000000000001"), -- i=4086
      ("11", "1010110001011101", "1010000010000001", "1010110011011101"), -- i=4087
      ("00", "1000101001001000", "0010110110100101", "1011011111101101"), -- i=4088
      ("01", "1000101001001000", "0010110110100101", "0101110010100011"), -- i=4089
      ("10", "1000101001001000", "0010110110100101", "0000100000000000"), -- i=4090
      ("11", "1000101001001000", "0010110110100101", "1010111111101101"), -- i=4091
      ("00", "1010000011000001", "1111011100000111", "1001011111001000"), -- i=4092
      ("01", "1010000011000001", "1111011100000111", "1010100110111010"), -- i=4093
      ("10", "1010000011000001", "1111011100000111", "1010000000000001"), -- i=4094
      ("11", "1010000011000001", "1111011100000111", "1111011111000111"), -- i=4095
      ("00", "0001100101000010", "0011001000110100", "0100101101110110"), -- i=4096
      ("01", "0001100101000010", "0011001000110100", "1110011100001110"), -- i=4097
      ("10", "0001100101000010", "0011001000110100", "0001000000000000"), -- i=4098
      ("11", "0001100101000010", "0011001000110100", "0011101101110110"), -- i=4099
      ("00", "1100010001001010", "1001111101010101", "0110001110011111"), -- i=4100
      ("01", "1100010001001010", "1001111101010101", "0010010011110101"), -- i=4101
      ("10", "1100010001001010", "1001111101010101", "1000010001000000"), -- i=4102
      ("11", "1100010001001010", "1001111101010101", "1101111101011111"), -- i=4103
      ("00", "0001101100111001", "1001010110101000", "1011000011100001"), -- i=4104
      ("01", "0001101100111001", "1001010110101000", "1000010110010001"), -- i=4105
      ("10", "0001101100111001", "1001010110101000", "0001000100101000"), -- i=4106
      ("11", "0001101100111001", "1001010110101000", "1001111110111001"), -- i=4107
      ("00", "1101111001010100", "0010001000110000", "0000000010000100"), -- i=4108
      ("01", "1101111001010100", "0010001000110000", "1011110000100100"), -- i=4109
      ("10", "1101111001010100", "0010001000110000", "0000001000010000"), -- i=4110
      ("11", "1101111001010100", "0010001000110000", "1111111001110100"), -- i=4111
      ("00", "0010110000011000", "0010000010011011", "0100110010110011"), -- i=4112
      ("01", "0010110000011000", "0010000010011011", "0000101101111101"), -- i=4113
      ("10", "0010110000011000", "0010000010011011", "0010000000011000"), -- i=4114
      ("11", "0010110000011000", "0010000010011011", "0010110010011011"), -- i=4115
      ("00", "0100010111110100", "1010010101011000", "1110101101001100"), -- i=4116
      ("01", "0100010111110100", "1010010101011000", "1010000010011100"), -- i=4117
      ("10", "0100010111110100", "1010010101011000", "0000010101010000"), -- i=4118
      ("11", "0100010111110100", "1010010101011000", "1110010111111100"), -- i=4119
      ("00", "1001001000011000", "1100000110100000", "0101001110111000"), -- i=4120
      ("01", "1001001000011000", "1100000110100000", "1101000001111000"), -- i=4121
      ("10", "1001001000011000", "1100000110100000", "1000000000000000"), -- i=4122
      ("11", "1001001000011000", "1100000110100000", "1101001110111000"), -- i=4123
      ("00", "1100010000000000", "0101101001000001", "0001111001000001"), -- i=4124
      ("01", "1100010000000000", "0101101001000001", "0110100110111111"), -- i=4125
      ("10", "1100010000000000", "0101101001000001", "0100000000000000"), -- i=4126
      ("11", "1100010000000000", "0101101001000001", "1101111001000001"), -- i=4127
      ("00", "1011101001001001", "1010011110010000", "0110000111011001"), -- i=4128
      ("01", "1011101001001001", "1010011110010000", "0001001010111001"), -- i=4129
      ("10", "1011101001001001", "1010011110010000", "1010001000000000"), -- i=4130
      ("11", "1011101001001001", "1010011110010000", "1011111111011001"), -- i=4131
      ("00", "0111001000110110", "1110001011101100", "0101010100100010"), -- i=4132
      ("01", "0111001000110110", "1110001011101100", "1000111101001010"), -- i=4133
      ("10", "0111001000110110", "1110001011101100", "0110001000100100"), -- i=4134
      ("11", "0111001000110110", "1110001011101100", "1111001011111110"), -- i=4135
      ("00", "0010010011001000", "0111110010010100", "1010000101011100"), -- i=4136
      ("01", "0010010011001000", "0111110010010100", "1010100000110100"), -- i=4137
      ("10", "0010010011001000", "0111110010010100", "0010010010000000"), -- i=4138
      ("11", "0010010011001000", "0111110010010100", "0111110011011100"), -- i=4139
      ("00", "1111111111010100", "1111110111010101", "1111110110101001"), -- i=4140
      ("01", "1111111111010100", "1111110111010101", "0000000111111111"), -- i=4141
      ("10", "1111111111010100", "1111110111010101", "1111110111010100"), -- i=4142
      ("11", "1111111111010100", "1111110111010101", "1111111111010101"), -- i=4143
      ("00", "0001010010001010", "1111011101011101", "0000101111100111"), -- i=4144
      ("01", "0001010010001010", "1111011101011101", "0001110100101101"), -- i=4145
      ("10", "0001010010001010", "1111011101011101", "0001010000001000"), -- i=4146
      ("11", "0001010010001010", "1111011101011101", "1111011111011111"), -- i=4147
      ("00", "1011010101000111", "0011110100011011", "1111001001100010"), -- i=4148
      ("01", "1011010101000111", "0011110100011011", "0111100000101100"), -- i=4149
      ("10", "1011010101000111", "0011110100011011", "0011010100000011"), -- i=4150
      ("11", "1011010101000111", "0011110100011011", "1011110101011111"), -- i=4151
      ("00", "0001101111111110", "0101111101110010", "0111101101110000"), -- i=4152
      ("01", "0001101111111110", "0101111101110010", "1011110010001100"), -- i=4153
      ("10", "0001101111111110", "0101111101110010", "0001101101110010"), -- i=4154
      ("11", "0001101111111110", "0101111101110010", "0101111111111110"), -- i=4155
      ("00", "0110100111000101", "0010100001000111", "1001001000001100"), -- i=4156
      ("01", "0110100111000101", "0010100001000111", "0100000101111110"), -- i=4157
      ("10", "0110100111000101", "0010100001000111", "0010100001000101"), -- i=4158
      ("11", "0110100111000101", "0010100001000111", "0110100111000111"), -- i=4159
      ("00", "1100110100000101", "1011000010000010", "0111110110000111"), -- i=4160
      ("01", "1100110100000101", "1011000010000010", "0001110010000011"), -- i=4161
      ("10", "1100110100000101", "1011000010000010", "1000000000000000"), -- i=4162
      ("11", "1100110100000101", "1011000010000010", "1111110110000111"), -- i=4163
      ("00", "0101111011101000", "1110101101101000", "0100101001010000"), -- i=4164
      ("01", "0101111011101000", "1110101101101000", "0111001110000000"), -- i=4165
      ("10", "0101111011101000", "1110101101101000", "0100101001101000"), -- i=4166
      ("11", "0101111011101000", "1110101101101000", "1111111111101000"), -- i=4167
      ("00", "0110011111101110", "1100000000011011", "0010100000001001"), -- i=4168
      ("01", "0110011111101110", "1100000000011011", "1010011111010011"), -- i=4169
      ("10", "0110011111101110", "1100000000011011", "0100000000001010"), -- i=4170
      ("11", "0110011111101110", "1100000000011011", "1110011111111111"), -- i=4171
      ("00", "1001111110101111", "1010000101011100", "0100000100001011"), -- i=4172
      ("01", "1001111110101111", "1010000101011100", "1111111001010011"), -- i=4173
      ("10", "1001111110101111", "1010000101011100", "1000000100001100"), -- i=4174
      ("11", "1001111110101111", "1010000101011100", "1011111111111111"), -- i=4175
      ("00", "0110001001111000", "0010100000111110", "1000101010110110"), -- i=4176
      ("01", "0110001001111000", "0010100000111110", "0011101000111010"), -- i=4177
      ("10", "0110001001111000", "0010100000111110", "0010000000111000"), -- i=4178
      ("11", "0110001001111000", "0010100000111110", "0110101001111110"), -- i=4179
      ("00", "0001000101110001", "0101101010001000", "0110101111111001"), -- i=4180
      ("01", "0001000101110001", "0101101010001000", "1011011011101001"), -- i=4181
      ("10", "0001000101110001", "0101101010001000", "0001000000000000"), -- i=4182
      ("11", "0001000101110001", "0101101010001000", "0101101111111001"), -- i=4183
      ("00", "0000010100010101", "1100000010100111", "1100010110111100"), -- i=4184
      ("01", "0000010100010101", "1100000010100111", "0100010001101110"), -- i=4185
      ("10", "0000010100010101", "1100000010100111", "0000000000000101"), -- i=4186
      ("11", "0000010100010101", "1100000010100111", "1100010110110111"), -- i=4187
      ("00", "1101111010101010", "0011110001010011", "0001101011111101"), -- i=4188
      ("01", "1101111010101010", "0011110001010011", "1010001001010111"), -- i=4189
      ("10", "1101111010101010", "0011110001010011", "0001110000000010"), -- i=4190
      ("11", "1101111010101010", "0011110001010011", "1111111011111011"), -- i=4191
      ("00", "0010100111100010", "0001111111001100", "0100100110101110"), -- i=4192
      ("01", "0010100111100010", "0001111111001100", "0000101000010110"), -- i=4193
      ("10", "0010100111100010", "0001111111001100", "0000100111000000"), -- i=4194
      ("11", "0010100111100010", "0001111111001100", "0011111111101110"), -- i=4195
      ("00", "0100010010101111", "0111100100010110", "1011110111000101"), -- i=4196
      ("01", "0100010010101111", "0111100100010110", "1100101110011001"), -- i=4197
      ("10", "0100010010101111", "0111100100010110", "0100000000000110"), -- i=4198
      ("11", "0100010010101111", "0111100100010110", "0111110110111111"), -- i=4199
      ("00", "0101111000010011", "1111001111011101", "0101000111110000"), -- i=4200
      ("01", "0101111000010011", "1111001111011101", "0110101000110110"), -- i=4201
      ("10", "0101111000010011", "1111001111011101", "0101001000010001"), -- i=4202
      ("11", "0101111000010011", "1111001111011101", "1111111111011111"), -- i=4203
      ("00", "0001011010101110", "0110101101110101", "1000001000100011"), -- i=4204
      ("01", "0001011010101110", "0110101101110101", "1010101100111001"), -- i=4205
      ("10", "0001011010101110", "0110101101110101", "0000001000100100"), -- i=4206
      ("11", "0001011010101110", "0110101101110101", "0111111111111111"), -- i=4207
      ("00", "0100001111001001", "0000001101010100", "0100011100011101"), -- i=4208
      ("01", "0100001111001001", "0000001101010100", "0100000001110101"), -- i=4209
      ("10", "0100001111001001", "0000001101010100", "0000001101000000"), -- i=4210
      ("11", "0100001111001001", "0000001101010100", "0100001111011101"), -- i=4211
      ("00", "0111100110001111", "1101001100110110", "0100110011000101"), -- i=4212
      ("01", "0111100110001111", "1101001100110110", "1010011001011001"), -- i=4213
      ("10", "0111100110001111", "1101001100110110", "0101000100000110"), -- i=4214
      ("11", "0111100110001111", "1101001100110110", "1111101110111111"), -- i=4215
      ("00", "0001011110010100", "0100101111011001", "0110001101101101"), -- i=4216
      ("01", "0001011110010100", "0100101111011001", "1100101110111011"), -- i=4217
      ("10", "0001011110010100", "0100101111011001", "0000001110010000"), -- i=4218
      ("11", "0001011110010100", "0100101111011001", "0101111111011101"), -- i=4219
      ("00", "0111010110001110", "0000110100010101", "1000001010100011"), -- i=4220
      ("01", "0111010110001110", "0000110100010101", "0110100001111001"), -- i=4221
      ("10", "0111010110001110", "0000110100010101", "0000010100000100"), -- i=4222
      ("11", "0111010110001110", "0000110100010101", "0111110110011111"), -- i=4223
      ("00", "1010101000001110", "0000010110001100", "1010111110011010"), -- i=4224
      ("01", "1010101000001110", "0000010110001100", "1010010010000010"), -- i=4225
      ("10", "1010101000001110", "0000010110001100", "0000000000001100"), -- i=4226
      ("11", "1010101000001110", "0000010110001100", "1010111110001110"), -- i=4227
      ("00", "1111101110101010", "0010001000110001", "0001110111011011"), -- i=4228
      ("01", "1111101110101010", "0010001000110001", "1101100101111001"), -- i=4229
      ("10", "1111101110101010", "0010001000110001", "0010001000100000"), -- i=4230
      ("11", "1111101110101010", "0010001000110001", "1111101110111011"), -- i=4231
      ("00", "1111001101010111", "0100011111101111", "0011101101000110"), -- i=4232
      ("01", "1111001101010111", "0100011111101111", "1010101101101000"), -- i=4233
      ("10", "1111001101010111", "0100011111101111", "0100001101000111"), -- i=4234
      ("11", "1111001101010111", "0100011111101111", "1111011111111111"), -- i=4235
      ("00", "1110011001001000", "1011011100000000", "1001110101001000"), -- i=4236
      ("01", "1110011001001000", "1011011100000000", "0010111101001000"), -- i=4237
      ("10", "1110011001001000", "1011011100000000", "1010011000000000"), -- i=4238
      ("11", "1110011001001000", "1011011100000000", "1111011101001000"), -- i=4239
      ("00", "1010001101011110", "1010110100010100", "0101000001110010"), -- i=4240
      ("01", "1010001101011110", "1010110100010100", "1111011001001010"), -- i=4241
      ("10", "1010001101011110", "1010110100010100", "1010000100010100"), -- i=4242
      ("11", "1010001101011110", "1010110100010100", "1010111101011110"), -- i=4243
      ("00", "0100110110011001", "0011010011111101", "1000001010010110"), -- i=4244
      ("01", "0100110110011001", "0011010011111101", "0001100010011100"), -- i=4245
      ("10", "0100110110011001", "0011010011111101", "0000010010011001"), -- i=4246
      ("11", "0100110110011001", "0011010011111101", "0111110111111101"), -- i=4247
      ("00", "1011011101000000", "1001011010111010", "0100110111111010"), -- i=4248
      ("01", "1011011101000000", "1001011010111010", "0010000010000110"), -- i=4249
      ("10", "1011011101000000", "1001011010111010", "1001011000000000"), -- i=4250
      ("11", "1011011101000000", "1001011010111010", "1011011111111010"), -- i=4251
      ("00", "0100000110101000", "0000010101100101", "0100011100001101"), -- i=4252
      ("01", "0100000110101000", "0000010101100101", "0011110001000011"), -- i=4253
      ("10", "0100000110101000", "0000010101100101", "0000000100100000"), -- i=4254
      ("11", "0100000110101000", "0000010101100101", "0100010111101101"), -- i=4255
      ("00", "0010100100101100", "1010100010000000", "1101000110101100"), -- i=4256
      ("01", "0010100100101100", "1010100010000000", "1000000010101100"), -- i=4257
      ("10", "0010100100101100", "1010100010000000", "0010100000000000"), -- i=4258
      ("11", "0010100100101100", "1010100010000000", "1010100110101100"), -- i=4259
      ("00", "1001110100100011", "0101011011000110", "1111001111101001"), -- i=4260
      ("01", "1001110100100011", "0101011011000110", "0100011001011101"), -- i=4261
      ("10", "1001110100100011", "0101011011000110", "0001010000000010"), -- i=4262
      ("11", "1001110100100011", "0101011011000110", "1101111111100111"), -- i=4263
      ("00", "0100010110000110", "1010000101100011", "1110011011101001"), -- i=4264
      ("01", "0100010110000110", "1010000101100011", "1010010000100011"), -- i=4265
      ("10", "0100010110000110", "1010000101100011", "0000000100000010"), -- i=4266
      ("11", "0100010110000110", "1010000101100011", "1110010111100111"), -- i=4267
      ("00", "0010110100111101", "1011001000110100", "1101111101110001"), -- i=4268
      ("01", "0010110100111101", "1011001000110100", "0111101100001001"), -- i=4269
      ("10", "0010110100111101", "1011001000110100", "0010000000110100"), -- i=4270
      ("11", "0010110100111101", "1011001000110100", "1011111100111101"), -- i=4271
      ("00", "0000110101001100", "1111111000011010", "0000101101100110"), -- i=4272
      ("01", "0000110101001100", "1111111000011010", "0000111100110010"), -- i=4273
      ("10", "0000110101001100", "1111111000011010", "0000110000001000"), -- i=4274
      ("11", "0000110101001100", "1111111000011010", "1111111101011110"), -- i=4275
      ("00", "1101110000111111", "1001100001011110", "0111010010011101"), -- i=4276
      ("01", "1101110000111111", "1001100001011110", "0100001111100001"), -- i=4277
      ("10", "1101110000111111", "1001100001011110", "1001100000011110"), -- i=4278
      ("11", "1101110000111111", "1001100001011110", "1101110001111111"), -- i=4279
      ("00", "0101001011101101", "1011010100011100", "0000100000001001"), -- i=4280
      ("01", "0101001011101101", "1011010100011100", "1001110111010001"), -- i=4281
      ("10", "0101001011101101", "1011010100011100", "0001000000001100"), -- i=4282
      ("11", "0101001011101101", "1011010100011100", "1111011111111101"), -- i=4283
      ("00", "1110010110100110", "0111100111100110", "0101111110001100"), -- i=4284
      ("01", "1110010110100110", "0111100111100110", "0110101111000000"), -- i=4285
      ("10", "1110010110100110", "0111100111100110", "0110000110100110"), -- i=4286
      ("11", "1110010110100110", "0111100111100110", "1111110111100110"), -- i=4287
      ("00", "1110110000010011", "1110110001010100", "1101100001100111"), -- i=4288
      ("01", "1110110000010011", "1110110001010100", "1111111110111111"), -- i=4289
      ("10", "1110110000010011", "1110110001010100", "1110110000010000"), -- i=4290
      ("11", "1110110000010011", "1110110001010100", "1110110001010111"), -- i=4291
      ("00", "0101101111100110", "1010000110100110", "1111110110001100"), -- i=4292
      ("01", "0101101111100110", "1010000110100110", "1011101001000000"), -- i=4293
      ("10", "0101101111100110", "1010000110100110", "0000000110100110"), -- i=4294
      ("11", "0101101111100110", "1010000110100110", "1111101111100110"), -- i=4295
      ("00", "0110100000011000", "1011111111001111", "0010011111100111"), -- i=4296
      ("01", "0110100000011000", "1011111111001111", "1010100001001001"), -- i=4297
      ("10", "0110100000011000", "1011111111001111", "0010100000001000"), -- i=4298
      ("11", "0110100000011000", "1011111111001111", "1111111111011111"), -- i=4299
      ("00", "0111000100101110", "0001001011001001", "1000001111110111"), -- i=4300
      ("01", "0111000100101110", "0001001011001001", "0101111001100101"), -- i=4301
      ("10", "0111000100101110", "0001001011001001", "0001000000001000"), -- i=4302
      ("11", "0111000100101110", "0001001011001001", "0111001111101111"), -- i=4303
      ("00", "0011100000011001", "0000111111110011", "0100100000001100"), -- i=4304
      ("01", "0011100000011001", "0000111111110011", "0010100000100110"), -- i=4305
      ("10", "0011100000011001", "0000111111110011", "0000100000010001"), -- i=4306
      ("11", "0011100000011001", "0000111111110011", "0011111111111011"), -- i=4307
      ("00", "0000010111000000", "1110111111101111", "1111010110101111"), -- i=4308
      ("01", "0000010111000000", "1110111111101111", "0001010111010001"), -- i=4309
      ("10", "0000010111000000", "1110111111101111", "0000010111000000"), -- i=4310
      ("11", "0000010111000000", "1110111111101111", "1110111111101111"), -- i=4311
      ("00", "0001101011110001", "1101010011111111", "1110111111110000"), -- i=4312
      ("01", "0001101011110001", "1101010011111111", "0100010111110010"), -- i=4313
      ("10", "0001101011110001", "1101010011111111", "0001000011110001"), -- i=4314
      ("11", "0001101011110001", "1101010011111111", "1101111011111111"), -- i=4315
      ("00", "1111011111000011", "1011101110110010", "1011001101110101"), -- i=4316
      ("01", "1111011111000011", "1011101110110010", "0011110000010001"), -- i=4317
      ("10", "1111011111000011", "1011101110110010", "1011001110000010"), -- i=4318
      ("11", "1111011111000011", "1011101110110010", "1111111111110011"), -- i=4319
      ("00", "1110110010000101", "1010010011101010", "1001000101101111"), -- i=4320
      ("01", "1110110010000101", "1010010011101010", "0100011110011011"), -- i=4321
      ("10", "1110110010000101", "1010010011101010", "1010010010000000"), -- i=4322
      ("11", "1110110010000101", "1010010011101010", "1110110011101111"), -- i=4323
      ("00", "1001000110011110", "1010011001001001", "0011011111100111"), -- i=4324
      ("01", "1001000110011110", "1010011001001001", "1110101101010101"), -- i=4325
      ("10", "1001000110011110", "1010011001001001", "1000000000001000"), -- i=4326
      ("11", "1001000110011110", "1010011001001001", "1011011111011111"), -- i=4327
      ("00", "1010110100100100", "1110111111011110", "1001110100000010"), -- i=4328
      ("01", "1010110100100100", "1110111111011110", "1011110101000110"), -- i=4329
      ("10", "1010110100100100", "1110111111011110", "1010110100000100"), -- i=4330
      ("11", "1010110100100100", "1110111111011110", "1110111111111110"), -- i=4331
      ("00", "0011110100111001", "0010011100100111", "0110010001100000"), -- i=4332
      ("01", "0011110100111001", "0010011100100111", "0001011000010010"), -- i=4333
      ("10", "0011110100111001", "0010011100100111", "0010010100100001"), -- i=4334
      ("11", "0011110100111001", "0010011100100111", "0011111100111111"), -- i=4335
      ("00", "1011001011110100", "1111011011101001", "1010100111011101"), -- i=4336
      ("01", "1011001011110100", "1111011011101001", "1011110000001011"), -- i=4337
      ("10", "1011001011110100", "1111011011101001", "1011001011100000"), -- i=4338
      ("11", "1011001011110100", "1111011011101001", "1111011011111101"), -- i=4339
      ("00", "0101001111001001", "0101010011000110", "1010100010001111"), -- i=4340
      ("01", "0101001111001001", "0101010011000110", "1111111100000011"), -- i=4341
      ("10", "0101001111001001", "0101010011000110", "0101000011000000"), -- i=4342
      ("11", "0101001111001001", "0101010011000110", "0101011111001111"), -- i=4343
      ("00", "0111110010100110", "1010011110011001", "0010010000111111"), -- i=4344
      ("01", "0111110010100110", "1010011110011001", "1101010100001101"), -- i=4345
      ("10", "0111110010100110", "1010011110011001", "0010010010000000"), -- i=4346
      ("11", "0111110010100110", "1010011110011001", "1111111110111111"), -- i=4347
      ("00", "0111101011100111", "1100100000000100", "0100001011101011"), -- i=4348
      ("01", "0111101011100111", "1100100000000100", "1011001011100011"), -- i=4349
      ("10", "0111101011100111", "1100100000000100", "0100100000000100"), -- i=4350
      ("11", "0111101011100111", "1100100000000100", "1111101011100111"), -- i=4351
      ("00", "1000100111101100", "0101011010100100", "1110000010010000"), -- i=4352
      ("01", "1000100111101100", "0101011010100100", "0011001101001000"), -- i=4353
      ("10", "1000100111101100", "0101011010100100", "0000000010100100"), -- i=4354
      ("11", "1000100111101100", "0101011010100100", "1101111111101100"), -- i=4355
      ("00", "1000000100101011", "0101101110111010", "1101110011100101"), -- i=4356
      ("01", "1000000100101011", "0101101110111010", "0010010101110001"), -- i=4357
      ("10", "1000000100101011", "0101101110111010", "0000000100101010"), -- i=4358
      ("11", "1000000100101011", "0101101110111010", "1101101110111011"), -- i=4359
      ("00", "1111001101100000", "1100101011010011", "1011111000110011"), -- i=4360
      ("01", "1111001101100000", "1100101011010011", "0010100010001101"), -- i=4361
      ("10", "1111001101100000", "1100101011010011", "1100001001000000"), -- i=4362
      ("11", "1111001101100000", "1100101011010011", "1111101111110011"), -- i=4363
      ("00", "0001010110010010", "1100010010001000", "1101101000011010"), -- i=4364
      ("01", "0001010110010010", "1100010010001000", "0101000100001010"), -- i=4365
      ("10", "0001010110010010", "1100010010001000", "0000010010000000"), -- i=4366
      ("11", "0001010110010010", "1100010010001000", "1101010110011010"), -- i=4367
      ("00", "0011100011101110", "0010100011001001", "0110000110110111"), -- i=4368
      ("01", "0011100011101110", "0010100011001001", "0001000000100101"), -- i=4369
      ("10", "0011100011101110", "0010100011001001", "0010100011001000"), -- i=4370
      ("11", "0011100011101110", "0010100011001001", "0011100011101111"), -- i=4371
      ("00", "0000011001000111", "1100111111100010", "1101011000101001"), -- i=4372
      ("01", "0000011001000111", "1100111111100010", "0011011001100101"), -- i=4373
      ("10", "0000011001000111", "1100111111100010", "0000011001000010"), -- i=4374
      ("11", "0000011001000111", "1100111111100010", "1100111111100111"), -- i=4375
      ("00", "1110001011011110", "0001011101011110", "1111101000111100"), -- i=4376
      ("01", "1110001011011110", "0001011101011110", "1100101110000000"), -- i=4377
      ("10", "1110001011011110", "0001011101011110", "0000001001011110"), -- i=4378
      ("11", "1110001011011110", "0001011101011110", "1111011111011110"), -- i=4379
      ("00", "1110110010111000", "0001010011100011", "0000000110011011"), -- i=4380
      ("01", "1110110010111000", "0001010011100011", "1101011111010101"), -- i=4381
      ("10", "1110110010111000", "0001010011100011", "0000010010100000"), -- i=4382
      ("11", "1110110010111000", "0001010011100011", "1111110011111011"), -- i=4383
      ("00", "0001111100010001", "1110001110101110", "0000001010111111"), -- i=4384
      ("01", "0001111100010001", "1110001110101110", "0011101101100011"), -- i=4385
      ("10", "0001111100010001", "1110001110101110", "0000001100000000"), -- i=4386
      ("11", "0001111100010001", "1110001110101110", "1111111110111111"), -- i=4387
      ("00", "0100111000000011", "0000010010000110", "0101001010001001"), -- i=4388
      ("01", "0100111000000011", "0000010010000110", "0100100101111101"), -- i=4389
      ("10", "0100111000000011", "0000010010000110", "0000010000000010"), -- i=4390
      ("11", "0100111000000011", "0000010010000110", "0100111010000111"), -- i=4391
      ("00", "0111100100011010", "1000001100011000", "1111110000110010"), -- i=4392
      ("01", "0111100100011010", "1000001100011000", "1111011000000010"), -- i=4393
      ("10", "0111100100011010", "1000001100011000", "0000000100011000"), -- i=4394
      ("11", "0111100100011010", "1000001100011000", "1111101100011010"), -- i=4395
      ("00", "0100000000011101", "1001001000101001", "1101001001000110"), -- i=4396
      ("01", "0100000000011101", "1001001000101001", "1010110111110100"), -- i=4397
      ("10", "0100000000011101", "1001001000101001", "0000000000001001"), -- i=4398
      ("11", "0100000000011101", "1001001000101001", "1101001000111101"), -- i=4399
      ("00", "0010100100110111", "0001000010110001", "0011100111101000"), -- i=4400
      ("01", "0010100100110111", "0001000010110001", "0001100010000110"), -- i=4401
      ("10", "0010100100110111", "0001000010110001", "0000000000110001"), -- i=4402
      ("11", "0010100100110111", "0001000010110001", "0011100110110111"), -- i=4403
      ("00", "1001010101001001", "0010000010010010", "1011010111011011"), -- i=4404
      ("01", "1001010101001001", "0010000010010010", "0111010010110111"), -- i=4405
      ("10", "1001010101001001", "0010000010010010", "0000000000000000"), -- i=4406
      ("11", "1001010101001001", "0010000010010010", "1011010111011011"), -- i=4407
      ("00", "0011101101011101", "1100101100001101", "0000011001101010"), -- i=4408
      ("01", "0011101101011101", "1100101100001101", "0111000001010000"), -- i=4409
      ("10", "0011101101011101", "1100101100001101", "0000101100001101"), -- i=4410
      ("11", "0011101101011101", "1100101100001101", "1111101101011101"), -- i=4411
      ("00", "0110100010111100", "1111101011001011", "0110001110000111"), -- i=4412
      ("01", "0110100010111100", "1111101011001011", "0110110111110001"), -- i=4413
      ("10", "0110100010111100", "1111101011001011", "0110100010001000"), -- i=4414
      ("11", "0110100010111100", "1111101011001011", "1111101011111111"), -- i=4415
      ("00", "1111110011010111", "1010011001001011", "1010001100100010"), -- i=4416
      ("01", "1111110011010111", "1010011001001011", "0101011010001100"), -- i=4417
      ("10", "1111110011010111", "1010011001001011", "1010010001000011"), -- i=4418
      ("11", "1111110011010111", "1010011001001011", "1111111011011111"), -- i=4419
      ("00", "1010100010000010", "0110001110011100", "0000110000011110"), -- i=4420
      ("01", "1010100010000010", "0110001110011100", "0100010011100110"), -- i=4421
      ("10", "1010100010000010", "0110001110011100", "0010000010000000"), -- i=4422
      ("11", "1010100010000010", "0110001110011100", "1110101110011110"), -- i=4423
      ("00", "1011010000101110", "0011110111000011", "1111000111110001"), -- i=4424
      ("01", "1011010000101110", "0011110111000011", "0111011001101011"), -- i=4425
      ("10", "1011010000101110", "0011110111000011", "0011010000000010"), -- i=4426
      ("11", "1011010000101110", "0011110111000011", "1011110111101111"), -- i=4427
      ("00", "1110001000000110", "0011000101110000", "0001001101110110"), -- i=4428
      ("01", "1110001000000110", "0011000101110000", "1011000010010110"), -- i=4429
      ("10", "1110001000000110", "0011000101110000", "0010000000000000"), -- i=4430
      ("11", "1110001000000110", "0011000101110000", "1111001101110110"), -- i=4431
      ("00", "1010010001010110", "0100111111011001", "1111010000101111"), -- i=4432
      ("01", "1010010001010110", "0100111111011001", "0101010001111101"), -- i=4433
      ("10", "1010010001010110", "0100111111011001", "0000010001010000"), -- i=4434
      ("11", "1010010001010110", "0100111111011001", "1110111111011111"), -- i=4435
      ("00", "0010011111010110", "1111111111100011", "0010011110111001"), -- i=4436
      ("01", "0010011111010110", "1111111111100011", "0010011111110011"), -- i=4437
      ("10", "0010011111010110", "1111111111100011", "0010011111000010"), -- i=4438
      ("11", "0010011111010110", "1111111111100011", "1111111111110111"), -- i=4439
      ("00", "1100000101011001", "1111010110111011", "1011011100010100"), -- i=4440
      ("01", "1100000101011001", "1111010110111011", "1100101110011110"), -- i=4441
      ("10", "1100000101011001", "1111010110111011", "1100000100011001"), -- i=4442
      ("11", "1100000101011001", "1111010110111011", "1111010111111011"), -- i=4443
      ("00", "0110000001110001", "0011101101010111", "1001101111001000"), -- i=4444
      ("01", "0110000001110001", "0011101101010111", "0010010100011010"), -- i=4445
      ("10", "0110000001110001", "0011101101010111", "0010000001010001"), -- i=4446
      ("11", "0110000001110001", "0011101101010111", "0111101101110111"), -- i=4447
      ("00", "0100100111111000", "0111100000011010", "1100001000010010"), -- i=4448
      ("01", "0100100111111000", "0111100000011010", "1101000111011110"), -- i=4449
      ("10", "0100100111111000", "0111100000011010", "0100100000011000"), -- i=4450
      ("11", "0100100111111000", "0111100000011010", "0111100111111010"), -- i=4451
      ("00", "1010111101001110", "1010111001000001", "0101110110001111"), -- i=4452
      ("01", "1010111101001110", "1010111001000001", "0000000100001101"), -- i=4453
      ("10", "1010111101001110", "1010111001000001", "1010111001000000"), -- i=4454
      ("11", "1010111101001110", "1010111001000001", "1010111101001111"), -- i=4455
      ("00", "1010111100000110", "1111100100100111", "1010100000101101"), -- i=4456
      ("01", "1010111100000110", "1111100100100111", "1011010111011111"), -- i=4457
      ("10", "1010111100000110", "1111100100100111", "1010100100000110"), -- i=4458
      ("11", "1010111100000110", "1111100100100111", "1111111100100111"), -- i=4459
      ("00", "1111001001100001", "1100001100011000", "1011010101111001"), -- i=4460
      ("01", "1111001001100001", "1100001100011000", "0010111101001001"), -- i=4461
      ("10", "1111001001100001", "1100001100011000", "1100001000000000"), -- i=4462
      ("11", "1111001001100001", "1100001100011000", "1111001101111001"), -- i=4463
      ("00", "1100111001100011", "0010101101011100", "1111100110111111"), -- i=4464
      ("01", "1100111001100011", "0010101101011100", "1010001100000111"), -- i=4465
      ("10", "1100111001100011", "0010101101011100", "0000101001000000"), -- i=4466
      ("11", "1100111001100011", "0010101101011100", "1110111101111111"), -- i=4467
      ("00", "0111111111000110", "0110000100001011", "1110000011010001"), -- i=4468
      ("01", "0111111111000110", "0110000100001011", "0001111010111011"), -- i=4469
      ("10", "0111111111000110", "0110000100001011", "0110000100000010"), -- i=4470
      ("11", "0111111111000110", "0110000100001011", "0111111111001111"), -- i=4471
      ("00", "1000110011101011", "1111001111011000", "1000000011000011"), -- i=4472
      ("01", "1000110011101011", "1111001111011000", "1001100100010011"), -- i=4473
      ("10", "1000110011101011", "1111001111011000", "1000000011001000"), -- i=4474
      ("11", "1000110011101011", "1111001111011000", "1111111111111011"), -- i=4475
      ("00", "0110100001100100", "0010010011101011", "1000110101001111"), -- i=4476
      ("01", "0110100001100100", "0010010011101011", "0100001101111001"), -- i=4477
      ("10", "0110100001100100", "0010010011101011", "0010000001100000"), -- i=4478
      ("11", "0110100001100100", "0010010011101011", "0110110011101111"), -- i=4479
      ("00", "0100011110111001", "0010011001100011", "0110111000011100"), -- i=4480
      ("01", "0100011110111001", "0010011001100011", "0010000101010110"), -- i=4481
      ("10", "0100011110111001", "0010011001100011", "0000011000100001"), -- i=4482
      ("11", "0100011110111001", "0010011001100011", "0110011111111011"), -- i=4483
      ("00", "1000010110101100", "1011101011110011", "0100000010011111"), -- i=4484
      ("01", "1000010110101100", "1011101011110011", "1100101010111001"), -- i=4485
      ("10", "1000010110101100", "1011101011110011", "1000000010100000"), -- i=4486
      ("11", "1000010110101100", "1011101011110011", "1011111111111111"), -- i=4487
      ("00", "0110101010001101", "1000000001010111", "1110101011100100"), -- i=4488
      ("01", "0110101010001101", "1000000001010111", "1110101000110110"), -- i=4489
      ("10", "0110101010001101", "1000000001010111", "0000000000000101"), -- i=4490
      ("11", "0110101010001101", "1000000001010111", "1110101011011111"), -- i=4491
      ("00", "1000000110111110", "0100100101011001", "1100101100010111"), -- i=4492
      ("01", "1000000110111110", "0100100101011001", "0011100001100101"), -- i=4493
      ("10", "1000000110111110", "0100100101011001", "0000000100011000"), -- i=4494
      ("11", "1000000110111110", "0100100101011001", "1100100111111111"), -- i=4495
      ("00", "1011011001000001", "1010011100000000", "0101110101000001"), -- i=4496
      ("01", "1011011001000001", "1010011100000000", "0000111101000001"), -- i=4497
      ("10", "1011011001000001", "1010011100000000", "1010011000000000"), -- i=4498
      ("11", "1011011001000001", "1010011100000000", "1011011101000001"), -- i=4499
      ("00", "1101101010011110", "0010111011001110", "0000100101101100"), -- i=4500
      ("01", "1101101010011110", "0010111011001110", "1010101111010000"), -- i=4501
      ("10", "1101101010011110", "0010111011001110", "0000101010001110"), -- i=4502
      ("11", "1101101010011110", "0010111011001110", "1111111011011110"), -- i=4503
      ("00", "0110011110010010", "0011010100111100", "1001110011001110"), -- i=4504
      ("01", "0110011110010010", "0011010100111100", "0011001001010110"), -- i=4505
      ("10", "0110011110010010", "0011010100111100", "0010010100010000"), -- i=4506
      ("11", "0110011110010010", "0011010100111100", "0111011110111110"), -- i=4507
      ("00", "1001101001001101", "1101001101100000", "0110110110101101"), -- i=4508
      ("01", "1001101001001101", "1101001101100000", "1100011011101101"), -- i=4509
      ("10", "1001101001001101", "1101001101100000", "1001001001000000"), -- i=4510
      ("11", "1001101001001101", "1101001101100000", "1101101101101101"), -- i=4511
      ("00", "0111101110101001", "1101001101100000", "0100111100001001"), -- i=4512
      ("01", "0111101110101001", "1101001101100000", "1010100001001001"), -- i=4513
      ("10", "0111101110101001", "1101001101100000", "0101001100100000"), -- i=4514
      ("11", "0111101110101001", "1101001101100000", "1111101111101001"), -- i=4515
      ("00", "0001111011010111", "1110110101011000", "0000110000101111"), -- i=4516
      ("01", "0001111011010111", "1110110101011000", "0011000101111111"), -- i=4517
      ("10", "0001111011010111", "1110110101011000", "0000110001010000"), -- i=4518
      ("11", "0001111011010111", "1110110101011000", "1111111111011111"), -- i=4519
      ("00", "1100010100110000", "1110101110110011", "1011000011100011"), -- i=4520
      ("01", "1100010100110000", "1110101110110011", "1101100101111101"), -- i=4521
      ("10", "1100010100110000", "1110101110110011", "1100000100110000"), -- i=4522
      ("11", "1100010100110000", "1110101110110011", "1110111110110011"), -- i=4523
      ("00", "1101011011000011", "0110011100010011", "0011110111010110"), -- i=4524
      ("01", "1101011011000011", "0110011100010011", "0110111110110000"), -- i=4525
      ("10", "1101011011000011", "0110011100010011", "0100011000000011"), -- i=4526
      ("11", "1101011011000011", "0110011100010011", "1111011111010011"), -- i=4527
      ("00", "0110000111011001", "1100110100000111", "0010111011100000"), -- i=4528
      ("01", "0110000111011001", "1100110100000111", "1001010011010010"), -- i=4529
      ("10", "0110000111011001", "1100110100000111", "0100000100000001"), -- i=4530
      ("11", "0110000111011001", "1100110100000111", "1110110111011111"), -- i=4531
      ("00", "0100011101101100", "0000010111101011", "0100110101010111"), -- i=4532
      ("01", "0100011101101100", "0000010111101011", "0100000110000001"), -- i=4533
      ("10", "0100011101101100", "0000010111101011", "0000010101101000"), -- i=4534
      ("11", "0100011101101100", "0000010111101011", "0100011111101111"), -- i=4535
      ("00", "0110010110100110", "1111010000110100", "0101100111011010"), -- i=4536
      ("01", "0110010110100110", "1111010000110100", "0111000101110010"), -- i=4537
      ("10", "0110010110100110", "1111010000110100", "0110010000100100"), -- i=4538
      ("11", "0110010110100110", "1111010000110100", "1111010110110110"), -- i=4539
      ("00", "0000110000101011", "0000110110101001", "0001100111010100"), -- i=4540
      ("01", "0000110000101011", "0000110110101001", "1111111010000010"), -- i=4541
      ("10", "0000110000101011", "0000110110101001", "0000110000101001"), -- i=4542
      ("11", "0000110000101011", "0000110110101001", "0000110110101011"), -- i=4543
      ("00", "0011111001011001", "1100010010001001", "0000001011100010"), -- i=4544
      ("01", "0011111001011001", "1100010010001001", "0111100111010000"), -- i=4545
      ("10", "0011111001011001", "1100010010001001", "0000010000001001"), -- i=4546
      ("11", "0011111001011001", "1100010010001001", "1111111011011001"), -- i=4547
      ("00", "1011111001100011", "0101111100100100", "0001110110000111"), -- i=4548
      ("01", "1011111001100011", "0101111100100100", "0101111100111111"), -- i=4549
      ("10", "1011111001100011", "0101111100100100", "0001111000100000"), -- i=4550
      ("11", "1011111001100011", "0101111100100100", "1111111101100111"), -- i=4551
      ("00", "0110011011010011", "0010111001110100", "1001010101000111"), -- i=4552
      ("01", "0110011011010011", "0010111001110100", "0011100001011111"), -- i=4553
      ("10", "0110011011010011", "0010111001110100", "0010011001010000"), -- i=4554
      ("11", "0110011011010011", "0010111001110100", "0110111011110111"), -- i=4555
      ("00", "1101111111001100", "1111101111111011", "1101101111000111"), -- i=4556
      ("01", "1101111111001100", "1111101111111011", "1110001111010001"), -- i=4557
      ("10", "1101111111001100", "1111101111111011", "1101101111001000"), -- i=4558
      ("11", "1101111111001100", "1111101111111011", "1111111111111111"), -- i=4559
      ("00", "0111111101010010", "1010001011110001", "0010001001000011"), -- i=4560
      ("01", "0111111101010010", "1010001011110001", "1101110001100001"), -- i=4561
      ("10", "0111111101010010", "1010001011110001", "0010001001010000"), -- i=4562
      ("11", "0111111101010010", "1010001011110001", "1111111111110011"), -- i=4563
      ("00", "1111000110011100", "0110110010000110", "0101111000100010"), -- i=4564
      ("01", "1111000110011100", "0110110010000110", "1000010100010110"), -- i=4565
      ("10", "1111000110011100", "0110110010000110", "0110000010000100"), -- i=4566
      ("11", "1111000110011100", "0110110010000110", "1111110110011110"), -- i=4567
      ("00", "1100010011010111", "0011100110000110", "1111111001011101"), -- i=4568
      ("01", "1100010011010111", "0011100110000110", "1000101101010001"), -- i=4569
      ("10", "1100010011010111", "0011100110000110", "0000000010000110"), -- i=4570
      ("11", "1100010011010111", "0011100110000110", "1111110111010111"), -- i=4571
      ("00", "1101110001011010", "0100000010000010", "0001110011011100"), -- i=4572
      ("01", "1101110001011010", "0100000010000010", "1001101111011000"), -- i=4573
      ("10", "1101110001011010", "0100000010000010", "0100000000000010"), -- i=4574
      ("11", "1101110001011010", "0100000010000010", "1101110011011010"), -- i=4575
      ("00", "0010111100010111", "0001110111011100", "0100110011110011"), -- i=4576
      ("01", "0010111100010111", "0001110111011100", "0001000100111011"), -- i=4577
      ("10", "0010111100010111", "0001110111011100", "0000110100010100"), -- i=4578
      ("11", "0010111100010111", "0001110111011100", "0011111111011111"), -- i=4579
      ("00", "1010110110001101", "1100011000000110", "0111001110010011"), -- i=4580
      ("01", "1010110110001101", "1100011000000110", "1110011110000111"), -- i=4581
      ("10", "1010110110001101", "1100011000000110", "1000010000000100"), -- i=4582
      ("11", "1010110110001101", "1100011000000110", "1110111110001111"), -- i=4583
      ("00", "0011000111001110", "0011000100110011", "0110001100000001"), -- i=4584
      ("01", "0011000111001110", "0011000100110011", "0000000010011011"), -- i=4585
      ("10", "0011000111001110", "0011000100110011", "0011000100000010"), -- i=4586
      ("11", "0011000111001110", "0011000100110011", "0011000111111111"), -- i=4587
      ("00", "0111100101111111", "0001110110111111", "1001011100111110"), -- i=4588
      ("01", "0111100101111111", "0001110110111111", "0101101111000000"), -- i=4589
      ("10", "0111100101111111", "0001110110111111", "0001100100111111"), -- i=4590
      ("11", "0111100101111111", "0001110110111111", "0111110111111111"), -- i=4591
      ("00", "0011101101001111", "0100101101001011", "1000011010011010"), -- i=4592
      ("01", "0011101101001111", "0100101101001011", "1111000000000100"), -- i=4593
      ("10", "0011101101001111", "0100101101001011", "0000101101001011"), -- i=4594
      ("11", "0011101101001111", "0100101101001011", "0111101101001111"), -- i=4595
      ("00", "1110000011010100", "0000011010010011", "1110011101100111"), -- i=4596
      ("01", "1110000011010100", "0000011010010011", "1101101001000001"), -- i=4597
      ("10", "1110000011010100", "0000011010010011", "0000000010010000"), -- i=4598
      ("11", "1110000011010100", "0000011010010011", "1110011011010111"), -- i=4599
      ("00", "1000111110100010", "1010110110000000", "0011110100100010"), -- i=4600
      ("01", "1000111110100010", "1010110110000000", "1110001000100010"), -- i=4601
      ("10", "1000111110100010", "1010110110000000", "1000110110000000"), -- i=4602
      ("11", "1000111110100010", "1010110110000000", "1010111110100010"), -- i=4603
      ("00", "0101001010110001", "0001011000011010", "0110100011001011"), -- i=4604
      ("01", "0101001010110001", "0001011000011010", "0011110010010111"), -- i=4605
      ("10", "0101001010110001", "0001011000011010", "0001001000010000"), -- i=4606
      ("11", "0101001010110001", "0001011000011010", "0101011010111011"), -- i=4607
      ("00", "0000110010100111", "0000101000100110", "0001011011001101"), -- i=4608
      ("01", "0000110010100111", "0000101000100110", "0000001010000001"), -- i=4609
      ("10", "0000110010100111", "0000101000100110", "0000100000100110"), -- i=4610
      ("11", "0000110010100111", "0000101000100110", "0000111010100111"), -- i=4611
      ("00", "1010010110011100", "1001011010001111", "0011110000101011"), -- i=4612
      ("01", "1010010110011100", "1001011010001111", "0000111100001101"), -- i=4613
      ("10", "1010010110011100", "1001011010001111", "1000010010001100"), -- i=4614
      ("11", "1010010110011100", "1001011010001111", "1011011110011111"), -- i=4615
      ("00", "1011100011100111", "1111100101110010", "1011001001011001"), -- i=4616
      ("01", "1011100011100111", "1111100101110010", "1011111101110101"), -- i=4617
      ("10", "1011100011100111", "1111100101110010", "1011100001100010"), -- i=4618
      ("11", "1011100011100111", "1111100101110010", "1111100111110111"), -- i=4619
      ("00", "0000101001101000", "1110111000110101", "1111100010011101"), -- i=4620
      ("01", "0000101001101000", "1110111000110101", "0001110000110011"), -- i=4621
      ("10", "0000101001101000", "1110111000110101", "0000101000100000"), -- i=4622
      ("11", "0000101001101000", "1110111000110101", "1110111001111101"), -- i=4623
      ("00", "1011110000100011", "1101010001110110", "1001000010011001"), -- i=4624
      ("01", "1011110000100011", "1101010001110110", "1110011110101101"), -- i=4625
      ("10", "1011110000100011", "1101010001110110", "1001010000100010"), -- i=4626
      ("11", "1011110000100011", "1101010001110110", "1111110001110111"), -- i=4627
      ("00", "1010110111010010", "0100011100111101", "1111010100001111"), -- i=4628
      ("01", "1010110111010010", "0100011100111101", "0110011010010101"), -- i=4629
      ("10", "1010110111010010", "0100011100111101", "0000010100010000"), -- i=4630
      ("11", "1010110111010010", "0100011100111101", "1110111111111111"), -- i=4631
      ("00", "1000010111010010", "1011010111111100", "0011101111001110"), -- i=4632
      ("01", "1000010111010010", "1011010111111100", "1100111111010110"), -- i=4633
      ("10", "1000010111010010", "1011010111111100", "1000010111010000"), -- i=4634
      ("11", "1000010111010010", "1011010111111100", "1011010111111110"), -- i=4635
      ("00", "1001011010011001", "0010101010110111", "1100000101010000"), -- i=4636
      ("01", "1001011010011001", "0010101010110111", "0110101111100010"), -- i=4637
      ("10", "1001011010011001", "0010101010110111", "0000001010010001"), -- i=4638
      ("11", "1001011010011001", "0010101010110111", "1011111010111111"), -- i=4639
      ("00", "0111001011111100", "1101000001001111", "0100001101001011"), -- i=4640
      ("01", "0111001011111100", "1101000001001111", "1010001010101101"), -- i=4641
      ("10", "0111001011111100", "1101000001001111", "0101000001001100"), -- i=4642
      ("11", "0111001011111100", "1101000001001111", "1111001011111111"), -- i=4643
      ("00", "0110111100111000", "1110010000100000", "0101001101011000"), -- i=4644
      ("01", "0110111100111000", "1110010000100000", "1000101100011000"), -- i=4645
      ("10", "0110111100111000", "1110010000100000", "0110010000100000"), -- i=4646
      ("11", "0110111100111000", "1110010000100000", "1110111100111000"), -- i=4647
      ("00", "0011101001000110", "0101111000101010", "1001100001110000"), -- i=4648
      ("01", "0011101001000110", "0101111000101010", "1101110000011100"), -- i=4649
      ("10", "0011101001000110", "0101111000101010", "0001101000000010"), -- i=4650
      ("11", "0011101001000110", "0101111000101010", "0111111001101110"), -- i=4651
      ("00", "1111001110010011", "1100111010000010", "1100001000010101"), -- i=4652
      ("01", "1111001110010011", "1100111010000010", "0010010100010001"), -- i=4653
      ("10", "1111001110010011", "1100111010000010", "1100001010000010"), -- i=4654
      ("11", "1111001110010011", "1100111010000010", "1111111110010011"), -- i=4655
      ("00", "1100001000010001", "0011010001110011", "1111011010000100"), -- i=4656
      ("01", "1100001000010001", "0011010001110011", "1000110110011110"), -- i=4657
      ("10", "1100001000010001", "0011010001110011", "0000000000010001"), -- i=4658
      ("11", "1100001000010001", "0011010001110011", "1111011001110011"), -- i=4659
      ("00", "1010110000111111", "0001111101010010", "1100101110010001"), -- i=4660
      ("01", "1010110000111111", "0001111101010010", "1000110011101101"), -- i=4661
      ("10", "1010110000111111", "0001111101010010", "0000110000010010"), -- i=4662
      ("11", "1010110000111111", "0001111101010010", "1011111101111111"), -- i=4663
      ("00", "1100100111110001", "0110000101110100", "0010101101100101"), -- i=4664
      ("01", "1100100111110001", "0110000101110100", "0110100001111101"), -- i=4665
      ("10", "1100100111110001", "0110000101110100", "0100000101110000"), -- i=4666
      ("11", "1100100111110001", "0110000101110100", "1110100111110101"), -- i=4667
      ("00", "0111101000101000", "0101111001101000", "1101100010010000"), -- i=4668
      ("01", "0111101000101000", "0101111001101000", "0001101111000000"), -- i=4669
      ("10", "0111101000101000", "0101111001101000", "0101101000101000"), -- i=4670
      ("11", "0111101000101000", "0101111001101000", "0111111001101000"), -- i=4671
      ("00", "1111110111110101", "0101010110100101", "0101001110011010"), -- i=4672
      ("01", "1111110111110101", "0101010110100101", "1010100001010000"), -- i=4673
      ("10", "1111110111110101", "0101010110100101", "0101010110100101"), -- i=4674
      ("11", "1111110111110101", "0101010110100101", "1111110111110101"), -- i=4675
      ("00", "0011011011000100", "0111110111001111", "1011010010010011"), -- i=4676
      ("01", "0011011011000100", "0111110111001111", "1011100011110101"), -- i=4677
      ("10", "0011011011000100", "0111110111001111", "0011010011000100"), -- i=4678
      ("11", "0011011011000100", "0111110111001111", "0111111111001111"), -- i=4679
      ("00", "1001111101111010", "1100100101010100", "0110100011001110"), -- i=4680
      ("01", "1001111101111010", "1100100101010100", "1101011000100110"), -- i=4681
      ("10", "1001111101111010", "1100100101010100", "1000100101010000"), -- i=4682
      ("11", "1001111101111010", "1100100101010100", "1101111101111110"), -- i=4683
      ("00", "0101011000101000", "0110111101000111", "1100010101101111"), -- i=4684
      ("01", "0101011000101000", "0110111101000111", "1110011011100001"), -- i=4685
      ("10", "0101011000101000", "0110111101000111", "0100011000000000"), -- i=4686
      ("11", "0101011000101000", "0110111101000111", "0111111101101111"), -- i=4687
      ("00", "1110110010000011", "1111000110101111", "1101111000110010"), -- i=4688
      ("01", "1110110010000011", "1111000110101111", "1111101011010100"), -- i=4689
      ("10", "1110110010000011", "1111000110101111", "1110000010000011"), -- i=4690
      ("11", "1110110010000011", "1111000110101111", "1111110110101111"), -- i=4691
      ("00", "0000100110001111", "0010100010101101", "0011001000111100"), -- i=4692
      ("01", "0000100110001111", "0010100010101101", "1110000011100010"), -- i=4693
      ("10", "0000100110001111", "0010100010101101", "0000100010001101"), -- i=4694
      ("11", "0000100110001111", "0010100010101101", "0010100110101111"), -- i=4695
      ("00", "1101001111001011", "1001111100000010", "0111001011001101"), -- i=4696
      ("01", "1101001111001011", "1001111100000010", "0011010011001001"), -- i=4697
      ("10", "1101001111001011", "1001111100000010", "1001001100000010"), -- i=4698
      ("11", "1101001111001011", "1001111100000010", "1101111111001011"), -- i=4699
      ("00", "1101101000111010", "0100001110101001", "0001110111100011"), -- i=4700
      ("01", "1101101000111010", "0100001110101001", "1001011010010001"), -- i=4701
      ("10", "1101101000111010", "0100001110101001", "0100001000101000"), -- i=4702
      ("11", "1101101000111010", "0100001110101001", "1101101110111011"), -- i=4703
      ("00", "0101000100010100", "1000110100100011", "1101111000110111"), -- i=4704
      ("01", "0101000100010100", "1000110100100011", "1100001111110001"), -- i=4705
      ("10", "0101000100010100", "1000110100100011", "0000000100000000"), -- i=4706
      ("11", "0101000100010100", "1000110100100011", "1101110100110111"), -- i=4707
      ("00", "0001010110111001", "1100100001010101", "1101111000001110"), -- i=4708
      ("01", "0001010110111001", "1100100001010101", "0100110101100100"), -- i=4709
      ("10", "0001010110111001", "1100100001010101", "0000000000010001"), -- i=4710
      ("11", "0001010110111001", "1100100001010101", "1101110111111101"), -- i=4711
      ("00", "0000001001101000", "1000011001101111", "1000100011010111"), -- i=4712
      ("01", "0000001001101000", "1000011001101111", "0111101111111001"), -- i=4713
      ("10", "0000001001101000", "1000011001101111", "0000001001101000"), -- i=4714
      ("11", "0000001001101000", "1000011001101111", "1000011001101111"), -- i=4715
      ("00", "1010111000000000", "0011110111000111", "1110101111000111"), -- i=4716
      ("01", "1010111000000000", "0011110111000111", "0111000000111001"), -- i=4717
      ("10", "1010111000000000", "0011110111000111", "0010110000000000"), -- i=4718
      ("11", "1010111000000000", "0011110111000111", "1011111111000111"), -- i=4719
      ("00", "0010010001000010", "1111100011000111", "0001110100001001"), -- i=4720
      ("01", "0010010001000010", "1111100011000111", "0010101101111011"), -- i=4721
      ("10", "0010010001000010", "1111100011000111", "0010000001000010"), -- i=4722
      ("11", "0010010001000010", "1111100011000111", "1111110011000111"), -- i=4723
      ("00", "0110000011010111", "1100111010100001", "0010111101111000"), -- i=4724
      ("01", "0110000011010111", "1100111010100001", "1001001000110110"), -- i=4725
      ("10", "0110000011010111", "1100111010100001", "0100000010000001"), -- i=4726
      ("11", "0110000011010111", "1100111010100001", "1110111011110111"), -- i=4727
      ("00", "0010011111100001", "0100001101101101", "0110101101001110"), -- i=4728
      ("01", "0010011111100001", "0100001101101101", "1110010001110100"), -- i=4729
      ("10", "0010011111100001", "0100001101101101", "0000001101100001"), -- i=4730
      ("11", "0010011111100001", "0100001101101101", "0110011111101101"), -- i=4731
      ("00", "0001001110001111", "0010101100010000", "0011111010011111"), -- i=4732
      ("01", "0001001110001111", "0010101100010000", "1110100001111111"), -- i=4733
      ("10", "0001001110001111", "0010101100010000", "0000001100000000"), -- i=4734
      ("11", "0001001110001111", "0010101100010000", "0011101110011111"), -- i=4735
      ("00", "1000010000111011", "0101001110111100", "1101011111110111"), -- i=4736
      ("01", "1000010000111011", "0101001110111100", "0011000001111111"), -- i=4737
      ("10", "1000010000111011", "0101001110111100", "0000000000111000"), -- i=4738
      ("11", "1000010000111011", "0101001110111100", "1101011110111111"), -- i=4739
      ("00", "0101000100000001", "1101010011111000", "0010010111111001"), -- i=4740
      ("01", "0101000100000001", "1101010011111000", "0111110000001001"), -- i=4741
      ("10", "0101000100000001", "1101010011111000", "0101000000000000"), -- i=4742
      ("11", "0101000100000001", "1101010011111000", "1101010111111001"), -- i=4743
      ("00", "0011011101001101", "0001111000001111", "0101010101011100"), -- i=4744
      ("01", "0011011101001101", "0001111000001111", "0001100100111110"), -- i=4745
      ("10", "0011011101001101", "0001111000001111", "0001011000001101"), -- i=4746
      ("11", "0011011101001101", "0001111000001111", "0011111101001111"), -- i=4747
      ("00", "1100000101000100", "1010111000010101", "0110111101011001"), -- i=4748
      ("01", "1100000101000100", "1010111000010101", "0001001100101111"), -- i=4749
      ("10", "1100000101000100", "1010111000010101", "1000000000000100"), -- i=4750
      ("11", "1100000101000100", "1010111000010101", "1110111101010101"), -- i=4751
      ("00", "1010101010110101", "0001111101010111", "1100101000001100"), -- i=4752
      ("01", "1010101010110101", "0001111101010111", "1000101101011110"), -- i=4753
      ("10", "1010101010110101", "0001111101010111", "0000101000010101"), -- i=4754
      ("11", "1010101010110101", "0001111101010111", "1011111111110111"), -- i=4755
      ("00", "0100001110101010", "1111001101011110", "0011011100001000"), -- i=4756
      ("01", "0100001110101010", "1111001101011110", "0101000001001100"), -- i=4757
      ("10", "0100001110101010", "1111001101011110", "0100001100001010"), -- i=4758
      ("11", "0100001110101010", "1111001101011110", "1111001111111110"), -- i=4759
      ("00", "0101001111100111", "0101101100111000", "1010111100011111"), -- i=4760
      ("01", "0101001111100111", "0101101100111000", "1111100010101111"), -- i=4761
      ("10", "0101001111100111", "0101101100111000", "0101001100100000"), -- i=4762
      ("11", "0101001111100111", "0101101100111000", "0101101111111111"), -- i=4763
      ("00", "0000110011100000", "0100101111110111", "0101100011010111"), -- i=4764
      ("01", "0000110011100000", "0100101111110111", "1100000011101001"), -- i=4765
      ("10", "0000110011100000", "0100101111110111", "0000100011100000"), -- i=4766
      ("11", "0000110011100000", "0100101111110111", "0100111111110111"), -- i=4767
      ("00", "0111010101100100", "0011100110101000", "1010111100001100"), -- i=4768
      ("01", "0111010101100100", "0011100110101000", "0011101110111100"), -- i=4769
      ("10", "0111010101100100", "0011100110101000", "0011000100100000"), -- i=4770
      ("11", "0111010101100100", "0011100110101000", "0111110111101100"), -- i=4771
      ("00", "1100110001001101", "0011010101110010", "0000000110111111"), -- i=4772
      ("01", "1100110001001101", "0011010101110010", "1001011011011011"), -- i=4773
      ("10", "1100110001001101", "0011010101110010", "0000010001000000"), -- i=4774
      ("11", "1100110001001101", "0011010101110010", "1111110101111111"), -- i=4775
      ("00", "1101101110110011", "0011111001100100", "0001101000010111"), -- i=4776
      ("01", "1101101110110011", "0011111001100100", "1001110101001111"), -- i=4777
      ("10", "1101101110110011", "0011111001100100", "0001101000100000"), -- i=4778
      ("11", "1101101110110011", "0011111001100100", "1111111111110111"), -- i=4779
      ("00", "0110010100000101", "1110001000111100", "0100011101000001"), -- i=4780
      ("01", "0110010100000101", "1110001000111100", "1000001011001001"), -- i=4781
      ("10", "0110010100000101", "1110001000111100", "0110000000000100"), -- i=4782
      ("11", "0110010100000101", "1110001000111100", "1110011100111101"), -- i=4783
      ("00", "0100111000010110", "1101001111000001", "0010000111010111"), -- i=4784
      ("01", "0100111000010110", "1101001111000001", "0111101001010101"), -- i=4785
      ("10", "0100111000010110", "1101001111000001", "0100001000000000"), -- i=4786
      ("11", "0100111000010110", "1101001111000001", "1101111111010111"), -- i=4787
      ("00", "0011011111110000", "1001001001100011", "1100101001010011"), -- i=4788
      ("01", "0011011111110000", "1001001001100011", "1010010110001101"), -- i=4789
      ("10", "0011011111110000", "1001001001100011", "0001001001100000"), -- i=4790
      ("11", "0011011111110000", "1001001001100011", "1011011111110011"), -- i=4791
      ("00", "1011000000111101", "0100100110100100", "1111100111100001"), -- i=4792
      ("01", "1011000000111101", "0100100110100100", "0110011010011001"), -- i=4793
      ("10", "1011000000111101", "0100100110100100", "0000000000100100"), -- i=4794
      ("11", "1011000000111101", "0100100110100100", "1111100110111101"), -- i=4795
      ("00", "0101010111111100", "1000101000100011", "1110000000011111"), -- i=4796
      ("01", "0101010111111100", "1000101000100011", "1100101111011001"), -- i=4797
      ("10", "0101010111111100", "1000101000100011", "0000000000100000"), -- i=4798
      ("11", "0101010111111100", "1000101000100011", "1101111111111111"), -- i=4799
      ("00", "0111111101011001", "1011100010101000", "0011100000000001"), -- i=4800
      ("01", "0111111101011001", "1011100010101000", "1100011010110001"), -- i=4801
      ("10", "0111111101011001", "1011100010101000", "0011100000001000"), -- i=4802
      ("11", "0111111101011001", "1011100010101000", "1111111111111001"), -- i=4803
      ("00", "0011001001110100", "0000110011011101", "0011111101010001"), -- i=4804
      ("01", "0011001001110100", "0000110011011101", "0010010110010111"), -- i=4805
      ("10", "0011001001110100", "0000110011011101", "0000000001010100"), -- i=4806
      ("11", "0011001001110100", "0000110011011101", "0011111011111101"), -- i=4807
      ("00", "0110101001101100", "1011000011000110", "0001101100110010"), -- i=4808
      ("01", "0110101001101100", "1011000011000110", "1011100110100110"), -- i=4809
      ("10", "0110101001101100", "1011000011000110", "0010000001000100"), -- i=4810
      ("11", "0110101001101100", "1011000011000110", "1111101011101110"), -- i=4811
      ("00", "1001011011010110", "0010111001100111", "1100010100111101"), -- i=4812
      ("01", "1001011011010110", "0010111001100111", "0110100001101111"), -- i=4813
      ("10", "1001011011010110", "0010111001100111", "0000011001000110"), -- i=4814
      ("11", "1001011011010110", "0010111001100111", "1011111011110111"), -- i=4815
      ("00", "0100001010110010", "0111100111111100", "1011110010101110"), -- i=4816
      ("01", "0100001010110010", "0111100111111100", "1100100010110110"), -- i=4817
      ("10", "0100001010110010", "0111100111111100", "0100000010110000"), -- i=4818
      ("11", "0100001010110010", "0111100111111100", "0111101111111110"), -- i=4819
      ("00", "1010101011000010", "1101111111100001", "1000101010100011"), -- i=4820
      ("01", "1010101011000010", "1101111111100001", "1100101011100001"), -- i=4821
      ("10", "1010101011000010", "1101111111100001", "1000101011000000"), -- i=4822
      ("11", "1010101011000010", "1101111111100001", "1111111111100011"), -- i=4823
      ("00", "0110011001101000", "0011010011000000", "1001101100101000"), -- i=4824
      ("01", "0110011001101000", "0011010011000000", "0011000110101000"), -- i=4825
      ("10", "0110011001101000", "0011010011000000", "0010010001000000"), -- i=4826
      ("11", "0110011001101000", "0011010011000000", "0111011011101000"), -- i=4827
      ("00", "1101101111011111", "0101100001110011", "0011010001010010"), -- i=4828
      ("01", "1101101111011111", "0101100001110011", "1000001101101100"), -- i=4829
      ("10", "1101101111011111", "0101100001110011", "0101100001010011"), -- i=4830
      ("11", "1101101111011111", "0101100001110011", "1101101111111111"), -- i=4831
      ("00", "0001010101110011", "0101011101010110", "0110110011001001"), -- i=4832
      ("01", "0001010101110011", "0101011101010110", "1011111000011101"), -- i=4833
      ("10", "0001010101110011", "0101011101010110", "0001010101010010"), -- i=4834
      ("11", "0001010101110011", "0101011101010110", "0101011101110111"), -- i=4835
      ("00", "0101001011001000", "1101110110011101", "0011000001100101"), -- i=4836
      ("01", "0101001011001000", "1101110110011101", "0111010100101011"), -- i=4837
      ("10", "0101001011001000", "1101110110011101", "0101000010001000"), -- i=4838
      ("11", "0101001011001000", "1101110110011101", "1101111111011101"), -- i=4839
      ("00", "1101010010010001", "1101110000111110", "1011000011001111"), -- i=4840
      ("01", "1101010010010001", "1101110000111110", "1111100001010011"), -- i=4841
      ("10", "1101010010010001", "1101110000111110", "1101010000010000"), -- i=4842
      ("11", "1101010010010001", "1101110000111110", "1101110010111111"), -- i=4843
      ("00", "0110101101100101", "1111101000010000", "0110010101110101"), -- i=4844
      ("01", "0110101101100101", "1111101000010000", "0111000101010101"), -- i=4845
      ("10", "0110101101100101", "1111101000010000", "0110101000000000"), -- i=4846
      ("11", "0110101101100101", "1111101000010000", "1111101101110101"), -- i=4847
      ("00", "0010000100011011", "1111010101010110", "0001011001110001"), -- i=4848
      ("01", "0010000100011011", "1111010101010110", "0010101111000101"), -- i=4849
      ("10", "0010000100011011", "1111010101010110", "0010000100010010"), -- i=4850
      ("11", "0010000100011011", "1111010101010110", "1111010101011111"), -- i=4851
      ("00", "0101100001000101", "0110010100101010", "1011110101101111"), -- i=4852
      ("01", "0101100001000101", "0110010100101010", "1111001100011011"), -- i=4853
      ("10", "0101100001000101", "0110010100101010", "0100000000000000"), -- i=4854
      ("11", "0101100001000101", "0110010100101010", "0111110101101111"), -- i=4855
      ("00", "0011110010001110", "0011111001110001", "0111101011111111"), -- i=4856
      ("01", "0011110010001110", "0011111001110001", "1111111000011101"), -- i=4857
      ("10", "0011110010001110", "0011111001110001", "0011110000000000"), -- i=4858
      ("11", "0011110010001110", "0011111001110001", "0011111011111111"), -- i=4859
      ("00", "1011000111010001", "0011100010000101", "1110101001010110"), -- i=4860
      ("01", "1011000111010001", "0011100010000101", "0111100101001100"), -- i=4861
      ("10", "1011000111010001", "0011100010000101", "0011000010000001"), -- i=4862
      ("11", "1011000111010001", "0011100010000101", "1011100111010101"), -- i=4863
      ("00", "1100010001010000", "0011100101101011", "1111110110111011"), -- i=4864
      ("01", "1100010001010000", "0011100101101011", "1000101011100101"), -- i=4865
      ("10", "1100010001010000", "0011100101101011", "0000000001000000"), -- i=4866
      ("11", "1100010001010000", "0011100101101011", "1111110101111011"), -- i=4867
      ("00", "0011001101110101", "1001010001001010", "1100011110111111"), -- i=4868
      ("01", "0011001101110101", "1001010001001010", "1001111100101011"), -- i=4869
      ("10", "0011001101110101", "1001010001001010", "0001000001000000"), -- i=4870
      ("11", "0011001101110101", "1001010001001010", "1011011101111111"), -- i=4871
      ("00", "0001111101110011", "0101010100001110", "0111010010000001"), -- i=4872
      ("01", "0001111101110011", "0101010100001110", "1100101001100101"), -- i=4873
      ("10", "0001111101110011", "0101010100001110", "0001010100000010"), -- i=4874
      ("11", "0001111101110011", "0101010100001110", "0101111101111111"), -- i=4875
      ("00", "0101001000011000", "0111111000100110", "1101000000111110"), -- i=4876
      ("01", "0101001000011000", "0111111000100110", "1101001111110010"), -- i=4877
      ("10", "0101001000011000", "0111111000100110", "0101001000000000"), -- i=4878
      ("11", "0101001000011000", "0111111000100110", "0111111000111110"), -- i=4879
      ("00", "1000100101101001", "1101111101000110", "0110100010101111"), -- i=4880
      ("01", "1000100101101001", "1101111101000110", "1010101000100011"), -- i=4881
      ("10", "1000100101101001", "1101111101000110", "1000100101000000"), -- i=4882
      ("11", "1000100101101001", "1101111101000110", "1101111101101111"), -- i=4883
      ("00", "1010100010000010", "1001101000010101", "0100001010010111"), -- i=4884
      ("01", "1010100010000010", "1001101000010101", "0000111001101101"), -- i=4885
      ("10", "1010100010000010", "1001101000010101", "1000100000000000"), -- i=4886
      ("11", "1010100010000010", "1001101000010101", "1011101010010111"), -- i=4887
      ("00", "1010010111101110", "0000101001111100", "1011000001101010"), -- i=4888
      ("01", "1010010111101110", "0000101001111100", "1001101101110010"), -- i=4889
      ("10", "1010010111101110", "0000101001111100", "0000000001101100"), -- i=4890
      ("11", "1010010111101110", "0000101001111100", "1010111111111110"), -- i=4891
      ("00", "0110111101111100", "0101011101100010", "1100011011011110"), -- i=4892
      ("01", "0110111101111100", "0101011101100010", "0001100000011010"), -- i=4893
      ("10", "0110111101111100", "0101011101100010", "0100011101100000"), -- i=4894
      ("11", "0110111101111100", "0101011101100010", "0111111101111110"), -- i=4895
      ("00", "0001011110001111", "1001110100001100", "1011010010011011"), -- i=4896
      ("01", "0001011110001111", "1001110100001100", "0111101010000011"), -- i=4897
      ("10", "0001011110001111", "1001110100001100", "0001010100001100"), -- i=4898
      ("11", "0001011110001111", "1001110100001100", "1001111110001111"), -- i=4899
      ("00", "0101100011010111", "0100111110011000", "1010100001101111"), -- i=4900
      ("01", "0101100011010111", "0100111110011000", "0000100100111111"), -- i=4901
      ("10", "0101100011010111", "0100111110011000", "0100100010010000"), -- i=4902
      ("11", "0101100011010111", "0100111110011000", "0101111111011111"), -- i=4903
      ("00", "1000011110011100", "1111100100111110", "1000000011011010"), -- i=4904
      ("01", "1000011110011100", "1111100100111110", "1000111001011110"), -- i=4905
      ("10", "1000011110011100", "1111100100111110", "1000000100011100"), -- i=4906
      ("11", "1000011110011100", "1111100100111110", "1111111110111110"), -- i=4907
      ("00", "0010110110100100", "1110000000111000", "0000110111011100"), -- i=4908
      ("01", "0010110110100100", "1110000000111000", "0100110101101100"), -- i=4909
      ("10", "0010110110100100", "1110000000111000", "0010000000100000"), -- i=4910
      ("11", "0010110110100100", "1110000000111000", "1110110110111100"), -- i=4911
      ("00", "1110101101110001", "1110101100110001", "1101011010100010"), -- i=4912
      ("01", "1110101101110001", "1110101100110001", "0000000001000000"), -- i=4913
      ("10", "1110101101110001", "1110101100110001", "1110101100110001"), -- i=4914
      ("11", "1110101101110001", "1110101100110001", "1110101101110001"), -- i=4915
      ("00", "1000000100111110", "0111101101101111", "1111110010101101"), -- i=4916
      ("01", "1000000100111110", "0111101101101111", "0000010111001111"), -- i=4917
      ("10", "1000000100111110", "0111101101101111", "0000000100101110"), -- i=4918
      ("11", "1000000100111110", "0111101101101111", "1111101101111111"), -- i=4919
      ("00", "1001100001011011", "0001000110001110", "1010100111101001"), -- i=4920
      ("01", "1001100001011011", "0001000110001110", "1000011011001101"), -- i=4921
      ("10", "1001100001011011", "0001000110001110", "0001000000001010"), -- i=4922
      ("11", "1001100001011011", "0001000110001110", "1001100111011111"), -- i=4923
      ("00", "1010010000000110", "1100011100101011", "0110101100110001"), -- i=4924
      ("01", "1010010000000110", "1100011100101011", "1101110011011011"), -- i=4925
      ("10", "1010010000000110", "1100011100101011", "1000010000000010"), -- i=4926
      ("11", "1010010000000110", "1100011100101011", "1110011100101111"), -- i=4927
      ("00", "1110010010001010", "1100010100010001", "1010100110011011"), -- i=4928
      ("01", "1110010010001010", "1100010100010001", "0001111101111001"), -- i=4929
      ("10", "1110010010001010", "1100010100010001", "1100010000000000"), -- i=4930
      ("11", "1110010010001010", "1100010100010001", "1110010110011011"), -- i=4931
      ("00", "1100000111010110", "0110010101000110", "0010011100011100"), -- i=4932
      ("01", "1100000111010110", "0110010101000110", "0101110010010000"), -- i=4933
      ("10", "1100000111010110", "0110010101000110", "0100000101000110"), -- i=4934
      ("11", "1100000111010110", "0110010101000110", "1110010111010110"), -- i=4935
      ("00", "1010100011000111", "0001101000100110", "1100001011101101"), -- i=4936
      ("01", "1010100011000111", "0001101000100110", "1000111010100001"), -- i=4937
      ("10", "1010100011000111", "0001101000100110", "0000100000000110"), -- i=4938
      ("11", "1010100011000111", "0001101000100110", "1011101011100111"), -- i=4939
      ("00", "1100000110100111", "0010101010100000", "1110110001000111"), -- i=4940
      ("01", "1100000110100111", "0010101010100000", "1001011100000111"), -- i=4941
      ("10", "1100000110100111", "0010101010100000", "0000000010100000"), -- i=4942
      ("11", "1100000110100111", "0010101010100000", "1110101110100111"), -- i=4943
      ("00", "1111001111111110", "1111011100110100", "1110101100110010"), -- i=4944
      ("01", "1111001111111110", "1111011100110100", "1111110011001010"), -- i=4945
      ("10", "1111001111111110", "1111011100110100", "1111001100110100"), -- i=4946
      ("11", "1111001111111110", "1111011100110100", "1111011111111110"), -- i=4947
      ("00", "0000110011011011", "1001111001100000", "1010101100111011"), -- i=4948
      ("01", "0000110011011011", "1001111001100000", "0110111001111011"), -- i=4949
      ("10", "0000110011011011", "1001111001100000", "0000110001000000"), -- i=4950
      ("11", "0000110011011011", "1001111001100000", "1001111011111011"), -- i=4951
      ("00", "1010011010110110", "0100000101001010", "1110100000000000"), -- i=4952
      ("01", "1010011010110110", "0100000101001010", "0110010101101100"), -- i=4953
      ("10", "1010011010110110", "0100000101001010", "0000000000000010"), -- i=4954
      ("11", "1010011010110110", "0100000101001010", "1110011111111110"), -- i=4955
      ("00", "1101111000101101", "1101010110111101", "1011001111101010"), -- i=4956
      ("01", "1101111000101101", "1101010110111101", "0000100001110000"), -- i=4957
      ("10", "1101111000101101", "1101010110111101", "1101010000101101"), -- i=4958
      ("11", "1101111000101101", "1101010110111101", "1101111110111101"), -- i=4959
      ("00", "0111101000001100", "1101000001010000", "0100101001011100"), -- i=4960
      ("01", "0111101000001100", "1101000001010000", "1010100110111100"), -- i=4961
      ("10", "0111101000001100", "1101000001010000", "0101000000000000"), -- i=4962
      ("11", "0111101000001100", "1101000001010000", "1111101001011100"), -- i=4963
      ("00", "0001100101000001", "0010010000000010", "0011110101000011"), -- i=4964
      ("01", "0001100101000001", "0010010000000010", "1111010100111111"), -- i=4965
      ("10", "0001100101000001", "0010010000000010", "0000000000000000"), -- i=4966
      ("11", "0001100101000001", "0010010000000010", "0011110101000011"), -- i=4967
      ("00", "0010101011011010", "0011001011110111", "0101110111010001"), -- i=4968
      ("01", "0010101011011010", "0011001011110111", "1111011111100011"), -- i=4969
      ("10", "0010101011011010", "0011001011110111", "0010001011010010"), -- i=4970
      ("11", "0010101011011010", "0011001011110111", "0011101011111111"), -- i=4971
      ("00", "1111010101000101", "1010000110101100", "1001011011110001"), -- i=4972
      ("01", "1111010101000101", "1010000110101100", "0101001110011001"), -- i=4973
      ("10", "1111010101000101", "1010000110101100", "1010000100000100"), -- i=4974
      ("11", "1111010101000101", "1010000110101100", "1111010111101101"), -- i=4975
      ("00", "0001111100001110", "0100100111110011", "0110100100000001"), -- i=4976
      ("01", "0001111100001110", "0100100111110011", "1101010100011011"), -- i=4977
      ("10", "0001111100001110", "0100100111110011", "0000100100000010"), -- i=4978
      ("11", "0001111100001110", "0100100111110011", "0101111111111111"), -- i=4979
      ("00", "1111011000101001", "0100000011011001", "0011011100000010"), -- i=4980
      ("01", "1111011000101001", "0100000011011001", "1011010101010000"), -- i=4981
      ("10", "1111011000101001", "0100000011011001", "0100000000001001"), -- i=4982
      ("11", "1111011000101001", "0100000011011001", "1111011011111001"), -- i=4983
      ("00", "1110000001101000", "0110100101010001", "0100100110111001"), -- i=4984
      ("01", "1110000001101000", "0110100101010001", "0111011100010111"), -- i=4985
      ("10", "1110000001101000", "0110100101010001", "0110000001000000"), -- i=4986
      ("11", "1110000001101000", "0110100101010001", "1110100101111001"), -- i=4987
      ("00", "1100100101100000", "0000000001100000", "1100100111000000"), -- i=4988
      ("01", "1100100101100000", "0000000001100000", "1100100100000000"), -- i=4989
      ("10", "1100100101100000", "0000000001100000", "0000000001100000"), -- i=4990
      ("11", "1100100101100000", "0000000001100000", "1100100101100000"), -- i=4991
      ("00", "0011010100010011", "1111110111101010", "0011001011111101"), -- i=4992
      ("01", "0011010100010011", "1111110111101010", "0011011100101001"), -- i=4993
      ("10", "0011010100010011", "1111110111101010", "0011010100000010"), -- i=4994
      ("11", "0011010100010011", "1111110111101010", "1111110111111011"), -- i=4995
      ("00", "1001110000100100", "1101001001010101", "0110111001111001"), -- i=4996
      ("01", "1001110000100100", "1101001001010101", "1100100111001111"), -- i=4997
      ("10", "1001110000100100", "1101001001010101", "1001000000000100"), -- i=4998
      ("11", "1001110000100100", "1101001001010101", "1101111001110101"), -- i=4999
      ("00", "0111001111011110", "1010110001000010", "0010000000100000"), -- i=5000
      ("01", "0111001111011110", "1010110001000010", "1100011110011100"), -- i=5001
      ("10", "0111001111011110", "1010110001000010", "0010000001000010"), -- i=5002
      ("11", "0111001111011110", "1010110001000010", "1111111111011110"), -- i=5003
      ("00", "0110101010111111", "1111010111000111", "0110000010000110"), -- i=5004
      ("01", "0110101010111111", "1111010111000111", "0111010011111000"), -- i=5005
      ("10", "0110101010111111", "1111010111000111", "0110000010000111"), -- i=5006
      ("11", "0110101010111111", "1111010111000111", "1111111111111111"), -- i=5007
      ("00", "1110111100001001", "0111110101011100", "0110110001100101"), -- i=5008
      ("01", "1110111100001001", "0111110101011100", "0111000110101101"), -- i=5009
      ("10", "1110111100001001", "0111110101011100", "0110110100001000"), -- i=5010
      ("11", "1110111100001001", "0111110101011100", "1111111101011101"), -- i=5011
      ("00", "1001100101001001", "1101011011111000", "0111000001000001"), -- i=5012
      ("01", "1001100101001001", "1101011011111000", "1100001001010001"), -- i=5013
      ("10", "1001100101001001", "1101011011111000", "1001000001001000"), -- i=5014
      ("11", "1001100101001001", "1101011011111000", "1101111111111001"), -- i=5015
      ("00", "1111010111011010", "1111010101001011", "1110101100100101"), -- i=5016
      ("01", "1111010111011010", "1111010101001011", "0000000010001111"), -- i=5017
      ("10", "1111010111011010", "1111010101001011", "1111010101001010"), -- i=5018
      ("11", "1111010111011010", "1111010101001011", "1111010111011011"), -- i=5019
      ("00", "1101111111011001", "0000010001101111", "1110010001001000"), -- i=5020
      ("01", "1101111111011001", "0000010001101111", "1101101101101010"), -- i=5021
      ("10", "1101111111011001", "0000010001101111", "0000010001001001"), -- i=5022
      ("11", "1101111111011001", "0000010001101111", "1101111111111111"));
  begin
    for i in patterns'range loop
      A <= patterns(i).A;
      B <= patterns(i).B;
      ALUOP <= patterns(i).ALUOP;
      wait for 10 ns;
      assert std_match(RESULT, patterns(i).RESULT) OR (RESULT = "ZZZZZZZZZZZZZZZZ" AND patterns(i).RESULT = "ZZZZZZZZZZZZZZZZ")
        report "wrong value for RESULT, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).RESULT) & ", found " & to_string(RESULT) severity error;assert std_match(FLAG, patterns(i).FLAG) OR (FLAG = "ZZZZ" AND patterns(i).FLAG = "ZZZZ")
        report "wrong value for FLAG, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).FLAG) & ", found " & to_string(FLAG) severity error;end loop;
    wait;
  end process;
end behav;
